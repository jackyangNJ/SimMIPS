module const_4(
	output [31:0]num
);

	assign num = 32'd4;

endmodule