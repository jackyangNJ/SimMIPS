module IM(
	input [31:0]if_pc_out,
	output [31:0]if_instr_out
);

	

endmodule