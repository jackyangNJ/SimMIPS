module SinglePortRam
(
	input clk_i,
	input we_i,
	input [11:0] adr_i, 
	input [3:0] be_i, 
	input [31:0] dat_i,
	output[31:0] dat_o
);
	
	// use a multi-dimensional packed array
	//to model individual bytes within the word
	// (* ram_init_file = "ram_init.mif" *) logic [3:0][7:0] ram[0:4095];
	logic [3:0][7:0] ram[0:4095];
	integer i;
	initial
	begin
		for(i=0;i<4096;i=i+1)
			ram[i] = 0;
ram[0]=32'h3c1d9f00; 
ram[1]=32'h27bd252c; 
ram[2]=32'h3c199f00; 
ram[3]=32'h27390258; 
ram[4]=32'h03200008; 
ram[5]=32'h00000000; 
ram[6]=32'h1000ffff; 
ram[7]=32'h00000000; 
ram[8]=32'h308400ff; 
ram[9]=32'h3c02b800; 
ram[10]=32'h904303fd; 
ram[11]=32'h30630020; 
ram[12]=32'h1060fffc; 
ram[13]=32'h00000000; 
ram[14]=32'ha04403f8; 
ram[15]=32'h03e00008; 
ram[16]=32'h00000000; 
ram[17]=32'h3c02b800; 
ram[18]=32'h2403ff80; 
ram[19]=32'ha04003f9; 
ram[20]=32'ha04303fb; 
ram[21]=32'h2403001b; 
ram[22]=32'ha04303f8; 
ram[23]=32'h24030003; 
ram[24]=32'ha04003f9; 
ram[25]=32'ha04303fb; 
ram[26]=32'h2403ffc7; 
ram[27]=32'ha04303fa; 
ram[28]=32'h2403000b; 
ram[29]=32'ha04303fc; 
ram[30]=32'h03e00008; 
ram[31]=32'h00000000; 
ram[32]=32'h90860000; 
ram[33]=32'h3c02b800; 
ram[34]=32'h10c0000a; 
ram[35]=32'h00000000; 
ram[36]=32'h904303fd; 
ram[37]=32'h30630020; 
ram[38]=32'h1060fffd; 
ram[39]=32'h00000000; 
ram[40]=32'ha04603f8; 
ram[41]=32'h24840001; 
ram[42]=32'h90860000; 
ram[43]=32'h14c0fff8; 
ram[44]=32'h00000000; 
ram[45]=32'h03e00008; 
ram[46]=32'h00000000; 
ram[47]=32'h27bdffe8; 
ram[48]=32'hafa60020; 
ram[49]=32'h3c069f00; 
ram[50]=32'hafa5001c; 
ram[51]=32'h24c60020; 
ram[52]=32'h27a5001c; 
ram[53]=32'hafbf0014; 
ram[54]=32'hafa70024; 
ram[55]=32'hafa40018; 
ram[56]=32'h0fc0048b; 
ram[57]=32'h00000000; 
ram[58]=32'h8fbf0014; 
ram[59]=32'h27bd0018; 
ram[60]=32'h03e00008; 
ram[61]=32'h00000000; 
ram[62]=32'h90020021; 
ram[63]=32'h304200ff; 
ram[64]=32'h03e00008; 
ram[65]=32'h00000000; 
ram[66]=32'h24020020; 
ram[67]=32'h2403000b; 
ram[68]=32'ha0430000; 
ram[69]=32'h90420000; 
ram[70]=32'h304200ff; 
ram[71]=32'h03e00008; 
ram[72]=32'h00000000; 
ram[73]=32'h24020020; 
ram[74]=32'h2403000a; 
ram[75]=32'ha0430000; 
ram[76]=32'h90420000; 
ram[77]=32'h304200ff; 
ram[78]=32'h03e00008; 
ram[79]=32'h00000000; 
ram[80]=32'h24020020; 
ram[81]=32'h2403000c; 
ram[82]=32'ha0430000; 
ram[83]=32'h90420000; 
ram[84]=32'h304200ff; 
ram[85]=32'h03e00008; 
ram[86]=32'h00000000; 
ram[87]=32'h240200a0; 
ram[88]=32'h2403000c; 
ram[89]=32'ha0430000; 
ram[90]=32'h90420000; 
ram[91]=32'h304200ff; 
ram[92]=32'h03e00008; 
ram[93]=32'h00000000; 
ram[94]=32'h40026000; 
ram[95]=32'h3442ff00; 
ram[96]=32'h40826000; 
ram[97]=32'h24030021; 
ram[98]=32'h240200a1; 
ram[99]=32'h240bffff; 
ram[100]=32'ha06b0000; 
ram[101]=32'h24060020; 
ram[102]=32'ha04b0000; 
ram[103]=32'h240400a0; 
ram[104]=32'h2405000a; 
ram[105]=32'h240a0011; 
ram[106]=32'h24090002; 
ram[107]=32'h24080003; 
ram[108]=32'h24070068; 
ram[109]=32'h240b0004; 
ram[110]=32'ha0ca0000; 
ram[111]=32'ha0690000; 
ram[112]=32'ha06b0000; 
ram[113]=32'ha0680000; 
ram[114]=32'ha08a0000; 
ram[115]=32'ha0450000; 
ram[116]=32'ha0490000; 
ram[117]=32'ha0480000; 
ram[118]=32'ha0c70000; 
ram[119]=32'ha0c50000; 
ram[120]=32'ha0870000; 
ram[121]=32'ha0850000; 
ram[122]=32'h03e00008; 
ram[123]=32'h00000000; 
ram[124]=32'h2403000c; 
ram[125]=32'ha0030020; 
ram[126]=32'h90020020; 
ram[127]=32'h24040002; 
ram[128]=32'h30420007; 
ram[129]=32'h1044000e; 
ram[130]=32'h00000000; 
ram[131]=32'h24030007; 
ram[132]=32'h14430009; 
ram[133]=32'h00000000; 
ram[134]=32'h2403000b; 
ram[135]=32'ha0030020; 
ram[136]=32'h90040020; 
ram[137]=32'h2403ffff; 
ram[138]=32'h00042600; 
ram[139]=32'h00042603; 
ram[140]=32'h28840000; 
ram[141]=32'h0064100a; 
ram[142]=32'h03e00008; 
ram[143]=32'h00000000; 
ram[144]=32'ha00300a0; 
ram[145]=32'h900200a0; 
ram[146]=32'h30420007; 
ram[147]=32'h24420008; 
ram[148]=32'h03e00008; 
ram[149]=32'h00000000; 
ram[150]=32'h27bdffe0; 
ram[151]=32'hafbf001c; 
ram[152]=32'hafb20018; 
ram[153]=32'hafb10014; 
ram[154]=32'hafb00010; 
ram[155]=32'h0fc00011; 
ram[156]=32'h00000000; 
ram[157]=32'h00001021; 
ram[158]=32'h40826000; 
ram[159]=32'h3c049f00; 
ram[160]=32'h248414e0; 
ram[161]=32'h0fc0002f; 
ram[162]=32'h00000000; 
ram[163]=32'h3c028400; 
ram[164]=32'h24440078; 
ram[165]=32'h304300ff; 
ram[166]=32'ha0430000; 
ram[167]=32'h24420001; 
ram[168]=32'h1444fffc; 
ram[169]=32'h00000000; 
ram[170]=32'h3c108400; 
ram[171]=32'h3c129f00; 
ram[172]=32'h265214f0; 
ram[173]=32'h26110078; 
ram[174]=32'h8e060000; 
ram[175]=32'h02002821; 
ram[176]=32'h02402021; 
ram[177]=32'h26100004; 
ram[178]=32'h0fc0002f; 
ram[179]=32'h00000000; 
ram[180]=32'h1611fff9; 
ram[181]=32'h00000000; 
ram[182]=32'h0bc000b6; 
ram[183]=32'h00000000; 
ram[184]=32'h27bdffe0; 
ram[185]=32'h3c04ffff; 
ram[186]=32'hafb20018; 
ram[187]=32'h3c129f00; 
ram[188]=32'hafb00010; 
ram[189]=32'hafbf001c; 
ram[190]=32'hafb10014; 
ram[191]=32'h00008021; 
ram[192]=32'h0fc000ec; 
ram[193]=32'h00000000; 
ram[194]=32'h26521500; 
ram[195]=32'h0bc000d0; 
ram[196]=32'h00000000; 
ram[197]=32'h0fc00008; 
ram[198]=32'h00000000; 
ram[199]=32'h2404000a; 
ram[200]=32'h0fc00008; 
ram[201]=32'h00000000; 
ram[202]=32'h26040010; 
ram[203]=32'h0fc000f2; 
ram[204]=32'h00000000; 
ram[205]=32'h26100001; 
ram[206]=32'h2a020010; 
ram[207]=32'h0002800a; 
ram[208]=32'h02002021; 
ram[209]=32'h0fc00103; 
ram[210]=32'h00000000; 
ram[211]=32'h02402021; 
ram[212]=32'h00408821; 
ram[213]=32'h0fc00020; 
ram[214]=32'h00000000; 
ram[215]=32'h26040030; 
ram[216]=32'h308400ff; 
ram[217]=32'h0fc00008; 
ram[218]=32'h00000000; 
ram[219]=32'h2404003d; 
ram[220]=32'h0fc00008; 
ram[221]=32'h00000000; 
ram[222]=32'h24040031; 
ram[223]=32'h1620ffe5; 
ram[224]=32'h00000000; 
ram[225]=32'h24040030; 
ram[226]=32'h0fc00008; 
ram[227]=32'h00000000; 
ram[228]=32'h2404000a; 
ram[229]=32'h0fc00008; 
ram[230]=32'h00000000; 
ram[231]=32'h26040010; 
ram[232]=32'h0fc000fa; 
ram[233]=32'h00000000; 
ram[234]=32'h0bc000cd; 
ram[235]=32'h00000000; 
ram[236]=32'h3c02b800; 
ram[237]=32'h2403ffff; 
ram[238]=32'hac440404; 
ram[239]=32'hac430400; 
ram[240]=32'h03e00008; 
ram[241]=32'h00000000; 
ram[242]=32'h3c02b800; 
ram[243]=32'h8c430400; 
ram[244]=32'h24050001; 
ram[245]=32'h00852004; 
ram[246]=32'h00831825; 
ram[247]=32'hac430400; 
ram[248]=32'h03e00008; 
ram[249]=32'h00000000; 
ram[250]=32'h3c02b800; 
ram[251]=32'h24050001; 
ram[252]=32'h8c430400; 
ram[253]=32'h00852004; 
ram[254]=32'h00042827; 
ram[255]=32'h00a31824; 
ram[256]=32'hac430400; 
ram[257]=32'h03e00008; 
ram[258]=32'h00000000; 
ram[259]=32'h3c02b800; 
ram[260]=32'h8c430400; 
ram[261]=32'h24020001; 
ram[262]=32'h00821004; 
ram[263]=32'h00431024; 
ram[264]=32'h03e00008; 
ram[265]=32'h00000000; 
ram[266]=32'h27bdffe8; 
ram[267]=32'hafbf0014; 
ram[268]=32'h40046800; 
ram[269]=32'h0004202b; 
ram[270]=32'h0fc00008; 
ram[271]=32'h00000000; 
ram[272]=32'h0fc00050; 
ram[273]=32'h00000000; 
ram[274]=32'h00402021; 
ram[275]=32'h0fc00008; 
ram[276]=32'h00000000; 
ram[277]=32'h90040060; 
ram[278]=32'h8fbf0014; 
ram[279]=32'h308400ff; 
ram[280]=32'h27bd0018; 
ram[281]=32'h0bc00008; 
ram[282]=32'h00000000; 
ram[283]=32'h3c039f00; 
ram[284]=32'h24630428; 
ram[285]=32'h00031900; 
ram[286]=32'h3c020800; 
ram[287]=32'h00031982; 
ram[288]=32'h00621825; 
ram[289]=32'h3c028000; 
ram[290]=32'hac430000; 
ram[291]=32'h03e00008; 
ram[292]=32'h00000000; 
ram[293]=32'h90820000; 
ram[294]=32'h10400009; 
ram[295]=32'h00000000; 
ram[296]=32'h00801021; 
ram[297]=32'h24420001; 
ram[298]=32'h90430000; 
ram[299]=32'h1460fffd; 
ram[300]=32'h00000000; 
ram[301]=32'h00441023; 
ram[302]=32'h03e00008; 
ram[303]=32'h00000000; 
ram[304]=32'h00001021; 
ram[305]=32'h03e00008; 
ram[306]=32'h00000000; 
ram[307]=32'h90a30000; 
ram[308]=32'h00801021; 
ram[309]=32'h00803021; 
ram[310]=32'h10600007; 
ram[311]=32'h00000000; 
ram[312]=32'h24c60001; 
ram[313]=32'h24a50001; 
ram[314]=32'ha0c3ffff; 
ram[315]=32'h90a30000; 
ram[316]=32'h1460fffb; 
ram[317]=32'h00000000; 
ram[318]=32'ha0c00000; 
ram[319]=32'h03e00008; 
ram[320]=32'h00000000; 
ram[321]=32'h90830000; 
ram[322]=32'h00801021; 
ram[323]=32'h10600014; 
ram[324]=32'h00000000; 
ram[325]=32'h00801821; 
ram[326]=32'h24630001; 
ram[327]=32'h90660000; 
ram[328]=32'h14c0fffd; 
ram[329]=32'h00000000; 
ram[330]=32'h00621823; 
ram[331]=32'h90a60000; 
ram[332]=32'h00431821; 
ram[333]=32'h10c00007; 
ram[334]=32'h00000000; 
ram[335]=32'h24630001; 
ram[336]=32'h24a50001; 
ram[337]=32'ha066ffff; 
ram[338]=32'h90a60000; 
ram[339]=32'h14c0fffb; 
ram[340]=32'h00000000; 
ram[341]=32'ha0600000; 
ram[342]=32'h03e00008; 
ram[343]=32'h00000000; 
ram[344]=32'h00001821; 
ram[345]=32'h0bc0014b; 
ram[346]=32'h00000000; 
ram[347]=32'h90a30000; 
ram[348]=32'h00801021; 
ram[349]=32'h10600012; 
ram[350]=32'h00000000; 
ram[351]=32'h18c00010; 
ram[352]=32'h00000000; 
ram[353]=32'h00a63021; 
ram[354]=32'h00803821; 
ram[355]=32'h0bc00167; 
ram[356]=32'h00000000; 
ram[357]=32'h10a60007; 
ram[358]=32'h00000000; 
ram[359]=32'h24e70001; 
ram[360]=32'h24a50001; 
ram[361]=32'ha0e3ffff; 
ram[362]=32'h90a30000; 
ram[363]=32'h1460fff9; 
ram[364]=32'h00000000; 
ram[365]=32'ha0e00000; 
ram[366]=32'h03e00008; 
ram[367]=32'h00000000; 
ram[368]=32'h00403821; 
ram[369]=32'h0bc0016d; 
ram[370]=32'h00000000; 
ram[371]=32'h90830000; 
ram[372]=32'h00801021; 
ram[373]=32'h1060001b; 
ram[374]=32'h00000000; 
ram[375]=32'h00801821; 
ram[376]=32'h24630001; 
ram[377]=32'h90670000; 
ram[378]=32'h14e0fffd; 
ram[379]=32'h00000000; 
ram[380]=32'h00621823; 
ram[381]=32'h90a70000; 
ram[382]=32'h00431821; 
ram[383]=32'h10e0000e; 
ram[384]=32'h00000000; 
ram[385]=32'h18c0000c; 
ram[386]=32'h00000000; 
ram[387]=32'h00a63021; 
ram[388]=32'h0bc00188; 
ram[389]=32'h00000000; 
ram[390]=32'h10a60007; 
ram[391]=32'h00000000; 
ram[392]=32'h24630001; 
ram[393]=32'h24a50001; 
ram[394]=32'ha067ffff; 
ram[395]=32'h90a70000; 
ram[396]=32'h14e0fff9; 
ram[397]=32'h00000000; 
ram[398]=32'ha0600000; 
ram[399]=32'h03e00008; 
ram[400]=32'h00000000; 
ram[401]=32'h00001821; 
ram[402]=32'h0bc0017d; 
ram[403]=32'h00000000; 
ram[404]=32'h0bc0019c; 
ram[405]=32'h00000000; 
ram[406]=32'h24a50001; 
ram[407]=32'h00c31023; 
ram[408]=32'h10600008; 
ram[409]=32'h00000000; 
ram[410]=32'h14400007; 
ram[411]=32'h00000000; 
ram[412]=32'h90860000; 
ram[413]=32'h90a30000; 
ram[414]=32'h24840001; 
ram[415]=32'h14c0fff6; 
ram[416]=32'h00000000; 
ram[417]=32'h00c31023; 
ram[418]=32'h03e00008; 
ram[419]=32'h00000000; 
ram[420]=32'h90830000; 
ram[421]=32'h1060001b; 
ram[422]=32'h00000000; 
ram[423]=32'h90a20000; 
ram[424]=32'h10400018; 
ram[425]=32'h00000000; 
ram[426]=32'h18c00016; 
ram[427]=32'h00000000; 
ram[428]=32'h00621023; 
ram[429]=32'h24840001; 
ram[430]=32'h24a50001; 
ram[431]=32'h1040000d; 
ram[432]=32'h00000000; 
ram[433]=32'h0bc001ca; 
ram[434]=32'h00000000; 
ram[435]=32'h90a70000; 
ram[436]=32'h24840001; 
ram[437]=32'h00671023; 
ram[438]=32'h10e0000a; 
ram[439]=32'h00000000; 
ram[440]=32'h10c0000e; 
ram[441]=32'h00000000; 
ram[442]=32'h24a50001; 
ram[443]=32'h1440000c; 
ram[444]=32'h00000000; 
ram[445]=32'h90830000; 
ram[446]=32'h24c6ffff; 
ram[447]=32'h1460fff3; 
ram[448]=32'h00000000; 
ram[449]=32'h10c00005; 
ram[450]=32'h00000000; 
ram[451]=32'h90a20000; 
ram[452]=32'h00621023; 
ram[453]=32'h03e00008; 
ram[454]=32'h00000000; 
ram[455]=32'h00001021; 
ram[456]=32'h03e00008; 
ram[457]=32'h00000000; 
ram[458]=32'h03e00008; 
ram[459]=32'h00000000; 
ram[460]=32'h00801021; 
ram[461]=32'h10c00009; 
ram[462]=32'h00000000; 
ram[463]=32'h00a63021; 
ram[464]=32'h00801821; 
ram[465]=32'h24a50001; 
ram[466]=32'h90a7ffff; 
ram[467]=32'h24630001; 
ram[468]=32'ha067ffff; 
ram[469]=32'h14a6fffb; 
ram[470]=32'h00000000; 
ram[471]=32'h03e00008; 
ram[472]=32'h00000000; 
ram[473]=32'h00801021; 
ram[474]=32'h24c7ffff; 
ram[475]=32'h00801821; 
ram[476]=32'h2408ffff; 
ram[477]=32'h10c00008; 
ram[478]=32'h00000000; 
ram[479]=32'h24a50004; 
ram[480]=32'h8ca6fffc; 
ram[481]=32'h24630004; 
ram[482]=32'h24e7ffff; 
ram[483]=32'hac66fffc; 
ram[484]=32'h14e8fffa; 
ram[485]=32'h00000000; 
ram[486]=32'h03e00008; 
ram[487]=32'h00000000; 
ram[488]=32'h00801021; 
ram[489]=32'h30a500ff; 
ram[490]=32'h10c00007; 
ram[491]=32'h00000000; 
ram[492]=32'h00863021; 
ram[493]=32'h00801821; 
ram[494]=32'h24630001; 
ram[495]=32'ha065ffff; 
ram[496]=32'h1466fffd; 
ram[497]=32'h00000000; 
ram[498]=32'h03e00008; 
ram[499]=32'h00000000; 
ram[500]=32'h00801021; 
ram[501]=32'h30a5ffff; 
ram[502]=32'h24c7ffff; 
ram[503]=32'h00801821; 
ram[504]=32'h2408ffff; 
ram[505]=32'h10c00006; 
ram[506]=32'h00000000; 
ram[507]=32'h24630002; 
ram[508]=32'h24e7ffff; 
ram[509]=32'ha465fffe; 
ram[510]=32'h14e8fffc; 
ram[511]=32'h00000000; 
ram[512]=32'h03e00008; 
ram[513]=32'h00000000; 
ram[514]=32'h18c00011; 
ram[515]=32'h00000000; 
ram[516]=32'h90870000; 
ram[517]=32'h90a20000; 
ram[518]=32'h00001821; 
ram[519]=32'h10e20007; 
ram[520]=32'h00000000; 
ram[521]=32'h0bc00217; 
ram[522]=32'h00000000; 
ram[523]=32'h90e70000; 
ram[524]=32'h90420000; 
ram[525]=32'h14e20009; 
ram[526]=32'h00000000; 
ram[527]=32'h24630001; 
ram[528]=32'h00833821; 
ram[529]=32'h00a31021; 
ram[530]=32'h1466fff8; 
ram[531]=32'h00000000; 
ram[532]=32'h00001021; 
ram[533]=32'h03e00008; 
ram[534]=32'h00000000; 
ram[535]=32'h00e21023; 
ram[536]=32'h03e00008; 
ram[537]=32'h00000000; 
ram[538]=32'haca00000; 
ram[539]=32'h90820000; 
ram[540]=32'h10400016; 
ram[541]=32'h00000000; 
ram[542]=32'h2443ffd0; 
ram[543]=32'h2c63000a; 
ram[544]=32'h10600015; 
ram[545]=32'h00000000; 
ram[546]=32'h00001821; 
ram[547]=32'h0bc00227; 
ram[548]=32'h00000000; 
ram[549]=32'h10c00010; 
ram[550]=32'h00000000; 
ram[551]=32'h00033040; 
ram[552]=32'h000318c0; 
ram[553]=32'h00c31821; 
ram[554]=32'h00621021; 
ram[555]=32'h2443ffd0; 
ram[556]=32'haca30000; 
ram[557]=32'h24840001; 
ram[558]=32'h90820000; 
ram[559]=32'h2446ffd0; 
ram[560]=32'h2cc6000a; 
ram[561]=32'h1440fff3; 
ram[562]=32'h00000000; 
ram[563]=32'h00001021; 
ram[564]=32'h03e00008; 
ram[565]=32'h00000000; 
ram[566]=32'h2402ffff; 
ram[567]=32'h03e00008; 
ram[568]=32'h00000000; 
ram[569]=32'h04800030; 
ram[570]=32'h00000000; 
ram[571]=32'h10800029; 
ram[572]=32'h00000000; 
ram[573]=32'h3c076666; 
ram[574]=32'h00801021; 
ram[575]=32'h00003021; 
ram[576]=32'h24e76667; 
ram[577]=32'h0bc00244; 
ram[578]=32'h00000000; 
ram[579]=32'h00603021; 
ram[580]=32'h00470018; 
ram[581]=32'h000217c3; 
ram[582]=32'h00001810; 
ram[583]=32'h00031883; 
ram[584]=32'h00621023; 
ram[585]=32'h24c30001; 
ram[586]=32'h1440fff8; 
ram[587]=32'h00000000; 
ram[588]=32'h00a62821; 
ram[589]=32'h3c096666; 
ram[590]=32'ha0a00001; 
ram[591]=32'h00a01021; 
ram[592]=32'h25296667; 
ram[593]=32'h00890018; 
ram[594]=32'h00043fc3; 
ram[595]=32'h00001810; 
ram[596]=32'h2442ffff; 
ram[597]=32'h00031883; 
ram[598]=32'h00671823; 
ram[599]=32'h000338c0; 
ram[600]=32'h00034040; 
ram[601]=32'h01074021; 
ram[602]=32'h24470001; 
ram[603]=32'h00882023; 
ram[604]=32'h00e63821; 
ram[605]=32'h24840030; 
ram[606]=32'h00e53823; 
ram[607]=32'ha0440001; 
ram[608]=32'h00602021; 
ram[609]=32'h1ce0ffef; 
ram[610]=32'h00000000; 
ram[611]=32'h03e00008; 
ram[612]=32'h00000000; 
ram[613]=32'h24020030; 
ram[614]=32'ha0a20000; 
ram[615]=32'ha0a00001; 
ram[616]=32'h03e00008; 
ram[617]=32'h00000000; 
ram[618]=32'h2402002d; 
ram[619]=32'ha0a20000; 
ram[620]=32'h00042023; 
ram[621]=32'h24a50001; 
ram[622]=32'h0bc0023d; 
ram[623]=32'h00000000; 
ram[624]=32'h27bdff98; 
ram[625]=32'hafb60058; 
ram[626]=32'h3c169f00; 
ram[627]=32'hafb7005c; 
ram[628]=32'hafb50054; 
ram[629]=32'hafb40050; 
ram[630]=32'hafb00040; 
ram[631]=32'hafbf0064; 
ram[632]=32'hafbe0060; 
ram[633]=32'hafb3004c; 
ram[634]=32'hafb20048; 
ram[635]=32'hafb10044; 
ram[636]=32'hafa40030; 
ram[637]=32'h00808021; 
ram[638]=32'h24150025; 
ram[639]=32'h24170063; 
ram[640]=32'h27b40010; 
ram[641]=32'h26d61518; 
ram[642]=32'h90a30000; 
ram[643]=32'h10600009; 
ram[644]=32'h00000000; 
ram[645]=32'h10750016; 
ram[646]=32'h00000000; 
ram[647]=32'ha2030000; 
ram[648]=32'h24a50001; 
ram[649]=32'h90a30000; 
ram[650]=32'h26100001; 
ram[651]=32'h1460fff9; 
ram[652]=32'h00000000; 
ram[653]=32'ha2000000; 
ram[654]=32'h8fa40030; 
ram[655]=32'h8fbf0064; 
ram[656]=32'h8fbe0060; 
ram[657]=32'h8fb7005c; 
ram[658]=32'h8fb60058; 
ram[659]=32'h8fb50054; 
ram[660]=32'h8fb40050; 
ram[661]=32'h8fb3004c; 
ram[662]=32'h8fb20048; 
ram[663]=32'h8fb10044; 
ram[664]=32'h8fb00040; 
ram[665]=32'h27bd0068; 
ram[666]=32'h0bc00125; 
ram[667]=32'h00000000; 
ram[668]=32'h90a20001; 
ram[669]=32'h24b10001; 
ram[670]=32'h00009821; 
ram[671]=32'h00009021; 
ram[672]=32'h00005821; 
ram[673]=32'h00005021; 
ram[674]=32'h0000f021; 
ram[675]=32'h240c0073; 
ram[676]=32'h24190075; 
ram[677]=32'h24180064; 
ram[678]=32'h240e006f; 
ram[679]=32'h2409002d; 
ram[680]=32'h24040001; 
ram[681]=32'h240d002e; 
ram[682]=32'h240f0030; 
ram[683]=32'h10570068; 
ram[684]=32'h00000000; 
ram[685]=32'h2c470064; 
ram[686]=32'h10e00010; 
ram[687]=32'h00000000; 
ram[688]=32'h10490085; 
ram[689]=32'h00000000; 
ram[690]=32'h2c47002e; 
ram[691]=32'h10e00057; 
ram[692]=32'h00000000; 
ram[693]=32'h10400072; 
ram[694]=32'h00000000; 
ram[695]=32'h145500ae; 
ram[696]=32'h00000000; 
ram[697]=32'h26220001; 
ram[698]=32'ha2150000; 
ram[699]=32'h00402821; 
ram[700]=32'h26100001; 
ram[701]=32'h0bc00282; 
ram[702]=32'h00000000; 
ram[703]=32'h104c007d; 
ram[704]=32'h00000000; 
ram[705]=32'h2c470074; 
ram[706]=32'h10e0009e; 
ram[707]=32'h00000000; 
ram[708]=32'h10580003; 
ram[709]=32'h00000000; 
ram[710]=32'h144e009f; 
ram[711]=32'h00000000; 
ram[712]=32'h8cc30000; 
ram[713]=32'h24c60004; 
ram[714]=32'h146000c6; 
ram[715]=32'h00000000; 
ram[716]=32'h24020030; 
ram[717]=32'ha3a20010; 
ram[718]=32'h24020001; 
ram[719]=32'h0053202a; 
ram[720]=32'h02603821; 
ram[721]=32'h00006021; 
ram[722]=32'h24030001; 
ram[723]=32'ha3a00011; 
ram[724]=32'h24050030; 
ram[725]=32'h24080001; 
ram[726]=32'h000b500b; 
ram[727]=32'h0044380a; 
ram[728]=32'h118300db; 
ram[729]=32'h00000000; 
ram[730]=32'h13c301ac; 
ram[731]=32'h00000000; 
ram[732]=32'h00f2182a; 
ram[733]=32'h10600193; 
ram[734]=32'h00000000; 
ram[735]=32'h02471823; 
ram[736]=32'h24040030; 
ram[737]=32'h24090020; 
ram[738]=32'h02031821; 
ram[739]=32'h012a200a; 
ram[740]=32'h26100001; 
ram[741]=32'ha204ffff; 
ram[742]=32'h1603fffd; 
ram[743]=32'h00000000; 
ram[744]=32'h0047202a; 
ram[745]=32'h10800170; 
ram[746]=32'h00000000; 
ram[747]=32'h00e28023; 
ram[748]=32'h00708021; 
ram[749]=32'h24020030; 
ram[750]=32'h24630001; 
ram[751]=32'ha062ffff; 
ram[752]=32'h1470fffd; 
ram[753]=32'h00000000; 
ram[754]=32'h02801021; 
ram[755]=32'h10a00005; 
ram[756]=32'h00000000; 
ram[757]=32'h24420001; 
ram[758]=32'h90430000; 
ram[759]=32'h1460fffd; 
ram[760]=32'h00000000; 
ram[761]=32'h02002021; 
ram[762]=32'h0bc002fd; 
ram[763]=32'h00000000; 
ram[764]=32'h00602021; 
ram[765]=32'h2442ffff; 
ram[766]=32'h90470000; 
ram[767]=32'h0282282b; 
ram[768]=32'h24830001; 
ram[769]=32'ha0870000; 
ram[770]=32'h14a0fff9; 
ram[771]=32'h00000000; 
ram[772]=32'h02088021; 
ram[773]=32'ha0800001; 
ram[774]=32'h26220001; 
ram[775]=32'ha2000000; 
ram[776]=32'h00402821; 
ram[777]=32'h0bc00282; 
ram[778]=32'h00000000; 
ram[779]=32'h104d006c; 
ram[780]=32'h00000000; 
ram[781]=32'h144f0058; 
ram[782]=32'h00000000; 
ram[783]=32'h92220001; 
ram[784]=32'h240a0001; 
ram[785]=32'h26310001; 
ram[786]=32'h1457ff9a; 
ram[787]=32'h00000000; 
ram[788]=32'h17c000b4; 
ram[789]=32'h00000000; 
ram[790]=32'h2a420002; 
ram[791]=32'h1440013f; 
ram[792]=32'h00000000; 
ram[793]=32'h2652ffff; 
ram[794]=32'h02129021; 
ram[795]=32'h24020020; 
ram[796]=32'h26100001; 
ram[797]=32'ha202ffff; 
ram[798]=32'h1612fffd; 
ram[799]=32'h00000000; 
ram[800]=32'h90c20000; 
ram[801]=32'h26500001; 
ram[802]=32'ha2420000; 
ram[803]=32'h26220001; 
ram[804]=32'h24c60004; 
ram[805]=32'h00402821; 
ram[806]=32'h0bc00282; 
ram[807]=32'h00000000; 
ram[808]=32'h8fbf0064; 
ram[809]=32'h8fbe0060; 
ram[810]=32'h8fb7005c; 
ram[811]=32'h8fb60058; 
ram[812]=32'h8fb50054; 
ram[813]=32'h8fb40050; 
ram[814]=32'h8fb3004c; 
ram[815]=32'h8fb20048; 
ram[816]=32'h8fb10044; 
ram[817]=32'h8fb00040; 
ram[818]=32'h00001021; 
ram[819]=32'h27bd0068; 
ram[820]=32'h03e00008; 
ram[821]=32'h00000000; 
ram[822]=32'h13c40126; 
ram[823]=32'h00000000; 
ram[824]=32'h92220001; 
ram[825]=32'h241e0001; 
ram[826]=32'h26310001; 
ram[827]=32'h0bc002ab; 
ram[828]=32'h00000000; 
ram[829]=32'h8cc50000; 
ram[830]=32'h24c60004; 
ram[831]=32'h00a02021; 
ram[832]=32'hafa60034; 
ram[833]=32'hafa50038; 
ram[834]=32'h0fc00125; 
ram[835]=32'h00000000; 
ram[836]=32'h00403021; 
ram[837]=32'h8fa50038; 
ram[838]=32'h12600003; 
ram[839]=32'h00000000; 
ram[840]=32'h0262102a; 
ram[841]=32'h0262300b; 
ram[842]=32'h17c000ab; 
ram[843]=32'h00000000; 
ram[844]=32'h00d2102a; 
ram[845]=32'h104000d8; 
ram[846]=32'h00000000; 
ram[847]=32'h02469023; 
ram[848]=32'h02129021; 
ram[849]=32'h24030020; 
ram[850]=32'h26100001; 
ram[851]=32'ha203ffff; 
ram[852]=32'h1612fffd; 
ram[853]=32'h00000000; 
ram[854]=32'h02402021; 
ram[855]=32'hafa60038; 
ram[856]=32'h0fc00133; 
ram[857]=32'h00000000; 
ram[858]=32'h8fa60038; 
ram[859]=32'h26220001; 
ram[860]=32'h02468021; 
ram[861]=32'h00402821; 
ram[862]=32'h8fa60034; 
ram[863]=32'h0bc00282; 
ram[864]=32'h00000000; 
ram[865]=32'h1059ff66; 
ram[866]=32'h00000000; 
ram[867]=32'h24070078; 
ram[868]=32'h1047ff63; 
ram[869]=32'h00000000; 
ram[870]=32'h2447ffd0; 
ram[871]=32'h30e200ff; 
ram[872]=32'h2c42000a; 
ram[873]=32'h104000f3; 
ram[874]=32'h00000000; 
ram[875]=32'h26310001; 
ram[876]=32'h00124040; 
ram[877]=32'h92220000; 
ram[878]=32'h001290c0; 
ram[879]=32'h01129021; 
ram[880]=32'h00f29021; 
ram[881]=32'h2447ffd0; 
ram[882]=32'h30e800ff; 
ram[883]=32'h2d08000a; 
ram[884]=32'h1500fff6; 
ram[885]=32'h00000000; 
ram[886]=32'h0bc002ab; 
ram[887]=32'h00000000; 
ram[888]=32'h116400e4; 
ram[889]=32'h00000000; 
ram[890]=32'h92220001; 
ram[891]=32'h10490061; 
ram[892]=32'h00000000; 
ram[893]=32'h2447ffd0; 
ram[894]=32'h30e800ff; 
ram[895]=32'h2d08000a; 
ram[896]=32'h26310001; 
ram[897]=32'h1100000c; 
ram[898]=32'h00000000; 
ram[899]=32'h26310001; 
ram[900]=32'h00134040; 
ram[901]=32'h92220000; 
ram[902]=32'h001398c0; 
ram[903]=32'h01139821; 
ram[904]=32'h00f39821; 
ram[905]=32'h2447ffd0; 
ram[906]=32'h30e800ff; 
ram[907]=32'h2d08000a; 
ram[908]=32'h1500fff6; 
ram[909]=32'h00000000; 
ram[910]=32'h240b0001; 
ram[911]=32'h0bc002ab; 
ram[912]=32'h00000000; 
ram[913]=32'h24040064; 
ram[914]=32'h10440059; 
ram[915]=32'h00000000; 
ram[916]=32'h24040075; 
ram[917]=32'h10440058; 
ram[918]=32'h00000000; 
ram[919]=32'h24040078; 
ram[920]=32'h10440072; 
ram[921]=32'h00000000; 
ram[922]=32'h3842006f; 
ram[923]=32'h24040008; 
ram[924]=32'h0002200b; 
ram[925]=32'h00006021; 
ram[926]=32'h00001021; 
ram[927]=32'h0064001b; 
ram[928]=32'h24420001; 
ram[929]=32'h02822821; 
ram[930]=32'h00003810; 
ram[931]=32'h00001812; 
ram[932]=32'h02c73821; 
ram[933]=32'h90e70000; 
ram[934]=32'ha0a7ffff; 
ram[935]=32'h1460fff7; 
ram[936]=32'h00000000; 
ram[937]=32'h00404021; 
ram[938]=32'h02821821; 
ram[939]=32'ha0600000; 
ram[940]=32'h0053202a; 
ram[941]=32'h02603821; 
ram[942]=32'h24030001; 
ram[943]=32'h93a50010; 
ram[944]=32'h000b500b; 
ram[945]=32'h0044380a; 
ram[946]=32'h1583ff27; 
ram[947]=32'h00000000; 
ram[948]=32'h24e90001; 
ram[949]=32'h13cc0073; 
ram[950]=32'h00000000; 
ram[951]=32'h114c0057; 
ram[952]=32'h00000000; 
ram[953]=32'h0132182a; 
ram[954]=32'h02002021; 
ram[955]=32'h10600008; 
ram[956]=32'h00000000; 
ram[957]=32'h02492023; 
ram[958]=32'h02042021; 
ram[959]=32'h24030020; 
ram[960]=32'h26100001; 
ram[961]=32'ha203ffff; 
ram[962]=32'h1604fffd; 
ram[963]=32'h00000000; 
ram[964]=32'h2409002d; 
ram[965]=32'h24830001; 
ram[966]=32'ha0890000; 
ram[967]=32'h0bc002e8; 
ram[968]=32'h00000000; 
ram[969]=32'h90c30000; 
ram[970]=32'h2a420002; 
ram[971]=32'h26040001; 
ram[972]=32'h24c60004; 
ram[973]=32'ha2030000; 
ram[974]=32'h144000aa; 
ram[975]=32'h00000000; 
ram[976]=32'h02128021; 
ram[977]=32'h00801021; 
ram[978]=32'h24030020; 
ram[979]=32'h24420001; 
ram[980]=32'ha043ffff; 
ram[981]=32'h1450fffd; 
ram[982]=32'h00000000; 
ram[983]=32'h2650ffff; 
ram[984]=32'h26220001; 
ram[985]=32'h00908021; 
ram[986]=32'h00402821; 
ram[987]=32'h0bc00282; 
ram[988]=32'h00000000; 
ram[989]=32'h92220002; 
ram[990]=32'h26310002; 
ram[991]=32'h2447ffd0; 
ram[992]=32'h2ce7000a; 
ram[993]=32'h10e0ffac; 
ram[994]=32'h00000000; 
ram[995]=32'h26310001; 
ram[996]=32'h92220000; 
ram[997]=32'h2447ffd0; 
ram[998]=32'h2ce7000a; 
ram[999]=32'h14e0fffb; 
ram[1000]=32'h00000000; 
ram[1001]=32'h240b0001; 
ram[1002]=32'h0bc002ab; 
ram[1003]=32'h00000000; 
ram[1004]=32'h04600035; 
ram[1005]=32'h00000000; 
ram[1006]=32'h00006021; 
ram[1007]=32'h2404000a; 
ram[1008]=32'h1460ffad; 
ram[1009]=32'h00000000; 
ram[1010]=32'h00004021; 
ram[1011]=32'h00001021; 
ram[1012]=32'h0bc003aa; 
ram[1013]=32'h00000000; 
ram[1014]=32'h02002021; 
ram[1015]=32'hafa60038; 
ram[1016]=32'h0fc00133; 
ram[1017]=32'h00000000; 
ram[1018]=32'h8fa60038; 
ram[1019]=32'h00d2182a; 
ram[1020]=32'h02061021; 
ram[1021]=32'h10600083; 
ram[1022]=32'h00000000; 
ram[1023]=32'h02463023; 
ram[1024]=32'h00468021; 
ram[1025]=32'h24030020; 
ram[1026]=32'h24420001; 
ram[1027]=32'ha043ffff; 
ram[1028]=32'h1450fffd; 
ram[1029]=32'h00000000; 
ram[1030]=32'h8fa60034; 
ram[1031]=32'h26220001; 
ram[1032]=32'h00402821; 
ram[1033]=32'h0bc00282; 
ram[1034]=32'h00000000; 
ram[1035]=32'h24040010; 
ram[1036]=32'h00006021; 
ram[1037]=32'h0bc0039e; 
ram[1038]=32'h00000000; 
ram[1039]=32'h240a002d; 
ram[1040]=32'h0132202a; 
ram[1041]=32'h26030001; 
ram[1042]=32'ha20a0000; 
ram[1043]=32'h1080fed4; 
ram[1044]=32'h00000000; 
ram[1045]=32'h26440001; 
ram[1046]=32'h00892023; 
ram[1047]=32'h02048021; 
ram[1048]=32'h240a0030; 
ram[1049]=32'h00602021; 
ram[1050]=32'h24840001; 
ram[1051]=32'ha08affff; 
ram[1052]=32'h1490fffd; 
ram[1053]=32'h00000000; 
ram[1054]=32'h02494823; 
ram[1055]=32'h00691821; 
ram[1056]=32'h0bc002e8; 
ram[1057]=32'h00000000; 
ram[1058]=32'h00031823; 
ram[1059]=32'h240c0001; 
ram[1060]=32'h0bc003ef; 
ram[1061]=32'h00000000; 
ram[1062]=32'h02009021; 
ram[1063]=32'h0bc00356; 
ram[1064]=32'h00000000; 
ram[1065]=32'h2407002d; 
ram[1066]=32'h26030001; 
ram[1067]=32'ha2070000; 
ram[1068]=32'h10800051; 
ram[1069]=32'h00000000; 
ram[1070]=32'h02621023; 
ram[1071]=32'h00625021; 
ram[1072]=32'h24020030; 
ram[1073]=32'h24630001; 
ram[1074]=32'ha062ffff; 
ram[1075]=32'h146afffd; 
ram[1076]=32'h00000000; 
ram[1077]=32'h02801021; 
ram[1078]=32'h10a00005; 
ram[1079]=32'h00000000; 
ram[1080]=32'h24420001; 
ram[1081]=32'h90430000; 
ram[1082]=32'h1460fffd; 
ram[1083]=32'h00000000; 
ram[1084]=32'h01402021; 
ram[1085]=32'h0bc00440; 
ram[1086]=32'h00000000; 
ram[1087]=32'h00602021; 
ram[1088]=32'h2442ffff; 
ram[1089]=32'h90470000; 
ram[1090]=32'h0282282b; 
ram[1091]=32'h24830001; 
ram[1092]=32'ha0870000; 
ram[1093]=32'h14a0fff9; 
ram[1094]=32'h00000000; 
ram[1095]=32'h0132182a; 
ram[1096]=32'ha0800001; 
ram[1097]=32'h01481021; 
ram[1098]=32'h10600029; 
ram[1099]=32'h00000000; 
ram[1100]=32'h02494823; 
ram[1101]=32'h00498021; 
ram[1102]=32'h24030020; 
ram[1103]=32'h24420001; 
ram[1104]=32'ha043ffff; 
ram[1105]=32'h1450fffd; 
ram[1106]=32'h00000000; 
ram[1107]=32'ha2000000; 
ram[1108]=32'h26220001; 
ram[1109]=32'h0bc00308; 
ram[1110]=32'h00000000; 
ram[1111]=32'h02009021; 
ram[1112]=32'h0bc00320; 
ram[1113]=32'h00000000; 
ram[1114]=32'h00608021; 
ram[1115]=32'h0bc002f2; 
ram[1116]=32'h00000000; 
ram[1117]=32'h0225102b; 
ram[1118]=32'h1440ffa8; 
ram[1119]=32'h00000000; 
ram[1120]=32'h26220001; 
ram[1121]=32'h02003821; 
ram[1122]=32'h00a02021; 
ram[1123]=32'h0bc00466; 
ram[1124]=32'h00000000; 
ram[1125]=32'h90830000; 
ram[1126]=32'h24e70001; 
ram[1127]=32'h24840001; 
ram[1128]=32'ha0e3ffff; 
ram[1129]=32'h1482fffb; 
ram[1130]=32'h00000000; 
ram[1131]=32'h02251823; 
ram[1132]=32'h24630001; 
ram[1133]=32'h02038021; 
ram[1134]=32'h00402821; 
ram[1135]=32'h0bc00282; 
ram[1136]=32'h00000000; 
ram[1137]=32'h02001821; 
ram[1138]=32'h0bc002e8; 
ram[1139]=32'h00000000; 
ram[1140]=32'h00408021; 
ram[1141]=32'ha2000000; 
ram[1142]=32'h26220001; 
ram[1143]=32'h0bc00308; 
ram[1144]=32'h00000000; 
ram[1145]=32'h26220001; 
ram[1146]=32'h00808021; 
ram[1147]=32'h00402821; 
ram[1148]=32'h0bc00282; 
ram[1149]=32'h00000000; 
ram[1150]=32'h00605021; 
ram[1151]=32'h0bc00435; 
ram[1152]=32'h00000000; 
ram[1153]=32'h00408021; 
ram[1154]=32'h26220001; 
ram[1155]=32'h8fa60034; 
ram[1156]=32'h00402821; 
ram[1157]=32'h0bc00282; 
ram[1158]=32'h00000000; 
ram[1159]=32'h00e04821; 
ram[1160]=32'h02001821; 
ram[1161]=32'h0bc0042c; 
ram[1162]=32'h00000000; 
ram[1163]=32'h27bdfbe0; 
ram[1164]=32'h00801821; 
ram[1165]=32'h00a01021; 
ram[1166]=32'h27a40010; 
ram[1167]=32'hafb10414; 
ram[1168]=32'h00602821; 
ram[1169]=32'h00c08821; 
ram[1170]=32'h00403021; 
ram[1171]=32'hafb20418; 
ram[1172]=32'hafb00410; 
ram[1173]=32'hafbf041c; 
ram[1174]=32'h0fc00270; 
ram[1175]=32'h00000000; 
ram[1176]=32'h93a40010; 
ram[1177]=32'h00409021; 
ram[1178]=32'h27b00010; 
ram[1179]=32'h10800007; 
ram[1180]=32'h00000000; 
ram[1181]=32'h26100001; 
ram[1182]=32'h0220f809; 
ram[1183]=32'h00000000; 
ram[1184]=32'h92040000; 
ram[1185]=32'h1480fffb; 
ram[1186]=32'h00000000; 
ram[1187]=32'h8fbf041c; 
ram[1188]=32'h02401021; 
ram[1189]=32'h8fb10414; 
ram[1190]=32'h8fb20418; 
ram[1191]=32'h8fb00410; 
ram[1192]=32'h27bd0420; 
ram[1193]=32'h03e00008; 
ram[1194]=32'h00000000; 
ram[1195]=32'h27bdffe8; 
ram[1196]=32'hafa60020; 
ram[1197]=32'h27a60020; 
ram[1198]=32'hafbf0014; 
ram[1199]=32'hafa70024; 
ram[1200]=32'hafa5001c; 
ram[1201]=32'h0fc00270; 
ram[1202]=32'h00000000; 
ram[1203]=32'h8fbf0014; 
ram[1204]=32'h27bd0018; 
ram[1205]=32'h03e00008; 
ram[1206]=32'h00000000; 
ram[1207]=32'h90a20000; 
ram[1208]=32'h10400018; 
ram[1209]=32'h00000000; 
ram[1210]=32'h00a01021; 
ram[1211]=32'h24420001; 
ram[1212]=32'h90430000; 
ram[1213]=32'h1460fffd; 
ram[1214]=32'h00000000; 
ram[1215]=32'h2442ffff; 
ram[1216]=32'h90470000; 
ram[1217]=32'h00a2302b; 
ram[1218]=32'h24830001; 
ram[1219]=32'ha0870000; 
ram[1220]=32'h10c00009; 
ram[1221]=32'h00000000; 
ram[1222]=32'h00602021; 
ram[1223]=32'h2442ffff; 
ram[1224]=32'h90470000; 
ram[1225]=32'h00a2302b; 
ram[1226]=32'h24830001; 
ram[1227]=32'ha0870000; 
ram[1228]=32'h14c0fff9; 
ram[1229]=32'h00000000; 
ram[1230]=32'ha0800001; 
ram[1231]=32'h03e00008; 
ram[1232]=32'h00000000; 
ram[1233]=32'h00a01021; 
ram[1234]=32'h0bc004c7; 
ram[1235]=32'h00000000; 
ram[1236]=32'h10800040; 
ram[1237]=32'h00000000; 
ram[1238]=32'h27bdffd0; 
ram[1239]=32'hafbf002c; 
ram[1240]=32'hafb10028; 
ram[1241]=32'hafb00024; 
ram[1242]=32'h04800036; 
ram[1243]=32'h00000000; 
ram[1244]=32'h00004821; 
ram[1245]=32'h3c056666; 
ram[1246]=32'h00003021; 
ram[1247]=32'h24a56667; 
ram[1248]=32'h0bc004e3; 
ram[1249]=32'h00000000; 
ram[1250]=32'h02003021; 
ram[1251]=32'h00850018; 
ram[1252]=32'h000417c3; 
ram[1253]=32'h00001810; 
ram[1254]=32'h00850018; 
ram[1255]=32'h00031883; 
ram[1256]=32'h00621823; 
ram[1257]=32'h00033840; 
ram[1258]=32'h00004010; 
ram[1259]=32'h000318c0; 
ram[1260]=32'h00e31821; 
ram[1261]=32'h00831823; 
ram[1262]=32'h24d00001; 
ram[1263]=32'h27a40010; 
ram[1264]=32'h00084083; 
ram[1265]=32'h00903821; 
ram[1266]=32'h24630030; 
ram[1267]=32'h01022023; 
ram[1268]=32'ha0e3ffff; 
ram[1269]=32'h1480ffec; 
ram[1270]=32'h00000000; 
ram[1271]=32'h15200012; 
ram[1272]=32'h00000000; 
ram[1273]=32'h2610ffff; 
ram[1274]=32'h2411ffff; 
ram[1275]=32'h27a40010; 
ram[1276]=32'h00901021; 
ram[1277]=32'h90440000; 
ram[1278]=32'h2610ffff; 
ram[1279]=32'h0fc00008; 
ram[1280]=32'h00000000; 
ram[1281]=32'h1611fff9; 
ram[1282]=32'h00000000; 
ram[1283]=32'h8fbf002c; 
ram[1284]=32'h8fb10028; 
ram[1285]=32'h8fb00024; 
ram[1286]=32'h2404000a; 
ram[1287]=32'h27bd0030; 
ram[1288]=32'h0bc00008; 
ram[1289]=32'h00000000; 
ram[1290]=32'h27a30010; 
ram[1291]=32'h00701021; 
ram[1292]=32'h2403002d; 
ram[1293]=32'h24d00002; 
ram[1294]=32'ha0430000; 
ram[1295]=32'h0bc004f9; 
ram[1296]=32'h00000000; 
ram[1297]=32'h00042023; 
ram[1298]=32'h24090001; 
ram[1299]=32'h0bc004dd; 
ram[1300]=32'h00000000; 
ram[1301]=32'h24040030; 
ram[1302]=32'h0bc00008; 
ram[1303]=32'h00000000; 
ram[1304]=32'h27bdffd8; 
ram[1305]=32'h27a20010; 
ram[1306]=32'h3c059f00; 
ram[1307]=32'h27a60018; 
ram[1308]=32'hafb10020; 
ram[1309]=32'hafbf0024; 
ram[1310]=32'hafb0001c; 
ram[1311]=32'h00408821; 
ram[1312]=32'h24a51508; 
ram[1313]=32'h3083000f; 
ram[1314]=32'h00a31821; 
ram[1315]=32'h90630000; 
ram[1316]=32'h24420001; 
ram[1317]=32'ha043ffff; 
ram[1318]=32'h00042102; 
ram[1319]=32'h1446fff9; 
ram[1320]=32'h00000000; 
ram[1321]=32'h27b00017; 
ram[1322]=32'h2631ffff; 
ram[1323]=32'h92040000; 
ram[1324]=32'h2610ffff; 
ram[1325]=32'h0fc00008; 
ram[1326]=32'h00000000; 
ram[1327]=32'h1611fffb; 
ram[1328]=32'h00000000; 
ram[1329]=32'h8fbf0024; 
ram[1330]=32'h8fb10020; 
ram[1331]=32'h8fb0001c; 
ram[1332]=32'h2404000a; 
ram[1333]=32'h27bd0028; 
ram[1334]=32'h0bc00008; 
ram[1335]=32'h00000000; 
ram[1336]=32'h6c6c6568; 
ram[1337]=32'h6f77206f; 
ram[1338]=32'h0a646c72; 
ram[1339]=32'h00000000; 
ram[1340]=32'h72646461; 
ram[1341]=32'h25783020; 
ram[1342]=32'h203d2078; 
ram[1343]=32'h000a7825; 
ram[1344]=32'h74726f70; 
ram[1345]=32'h00000000; 
ram[1346]=32'h33323130; 
ram[1347]=32'h37363534; 
ram[1348]=32'h62613938; 
ram[1349]=32'h66656463; 
ram[1350]=32'h33323130; 
ram[1351]=32'h37363534; 
ram[1352]=32'h42413938; 
ram[1353]=32'h46454443; 
ram[1354]=32'h00000000; 


	end
	
	reg[31:0] q;
	always_ff@(posedge clk_i)
	begin
	if(we_i) 
		begin
			if(be_i[0]) ram[adr_i][0] <= dat_i[7:0];
			if(be_i[1]) ram[adr_i][1] <= dat_i[15:8];
			if(be_i[2]) ram[adr_i][2] <= dat_i[23:16];
			if(be_i[3]) ram[adr_i][3] <= dat_i[31:24];
		end
		q <= ram[adr_i];
	end
	
	assign dat_o = q;
endmodule
