module DM(
	input mem_dmen,
	input mem_memwr,
	input [31:0]mem_result,
	input [31:0]mem_rt,
	output [31:0]mem_dout
);

endmodule