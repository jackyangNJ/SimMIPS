module const_base(
	output [31:0]base
);

	assign base = 32'h8000_0000;

endmodule