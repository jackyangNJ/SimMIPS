module SinglePortRam
(
	input clk_i,
	input we_i,
	input [11:0] adr_i, 
	input [3:0] be_i, 
	input [31:0] dat_i,
	output[31:0] dat_o
);
	
	// use a multi-dimensional packed array
	//to model individual bytes within the word
	// (* ram_init_file = "ram_init.mif" *) logic [3:0][7:0] ram[0:4095];
	logic [3:0][7:0] ram[0:4095];
	integer i;
	initial
	begin
		for(i=0;i<4096;i=i+1)
			ram[i] = 0;
			ram[0]=32'h3c1d9f00; 
ram[0]=32'h3c1d9f00; 
ram[1]=32'h27bd3fe8; 
ram[2]=32'h3c199f00; 
ram[3]=32'h27390198; 
ram[4]=32'h03200008; 
ram[5]=32'h00000000; 
ram[6]=32'h1000ffff; 
ram[7]=32'h00000000; 
ram[8]=32'h27bdffe0; 
ram[9]=32'h24020001; 
ram[10]=32'hafbf001c; 
ram[11]=32'hafb20018; 
ram[12]=32'hafb10014; 
ram[13]=32'hafb00010; 
ram[14]=32'h10c2000e; 
ram[15]=32'h00000000; 
ram[16]=32'h24020002; 
ram[17]=32'h10c20021; 
ram[18]=32'h00000000; 
ram[19]=32'h24020004; 
ram[20]=32'h10c20038; 
ram[21]=32'h00000000; 
ram[22]=32'h8fbf001c; 
ram[23]=32'h8fb20018; 
ram[24]=32'h8fb10014; 
ram[25]=32'h8fb00010; 
ram[26]=32'h27bd0020; 
ram[27]=32'h03e00008; 
ram[28]=32'h00000000; 
ram[29]=32'h18a0fff8; 
ram[30]=32'h00000000; 
ram[31]=32'h3c119f00; 
ram[32]=32'h00a49021; 
ram[33]=32'h00808021; 
ram[34]=32'h263128a0; 
ram[35]=32'h92060000; 
ram[36]=32'h02002821; 
ram[37]=32'h02202021; 
ram[38]=32'h26100001; 
ram[39]=32'h30c600ff; 
ram[40]=32'h0fc00254; 
ram[41]=32'h00000000; 
ram[42]=32'h1612fff8; 
ram[43]=32'h00000000; 
ram[44]=32'h8fbf001c; 
ram[45]=32'h8fb20018; 
ram[46]=32'h8fb10014; 
ram[47]=32'h8fb00010; 
ram[48]=32'h27bd0020; 
ram[49]=32'h03e00008; 
ram[50]=32'h00000000; 
ram[51]=32'h18a0ffe2; 
ram[52]=32'h00000000; 
ram[53]=32'h24a2ffff; 
ram[54]=32'h00021042; 
ram[55]=32'h24920002; 
ram[56]=32'h00021040; 
ram[57]=32'h3c119f00; 
ram[58]=32'h02429021; 
ram[59]=32'h00808021; 
ram[60]=32'h263128a0; 
ram[61]=32'h96060000; 
ram[62]=32'h02002821; 
ram[63]=32'h02202021; 
ram[64]=32'h26100002; 
ram[65]=32'h30c6ffff; 
ram[66]=32'h0fc00254; 
ram[67]=32'h00000000; 
ram[68]=32'h1612fff8; 
ram[69]=32'h00000000; 
ram[70]=32'h8fbf001c; 
ram[71]=32'h8fb20018; 
ram[72]=32'h8fb10014; 
ram[73]=32'h8fb00010; 
ram[74]=32'h27bd0020; 
ram[75]=32'h03e00008; 
ram[76]=32'h00000000; 
ram[77]=32'h18a0ffc8; 
ram[78]=32'h00000000; 
ram[79]=32'h24a2ffff; 
ram[80]=32'h00021082; 
ram[81]=32'h24920004; 
ram[82]=32'h00021080; 
ram[83]=32'h3c119f00; 
ram[84]=32'h02429021; 
ram[85]=32'h00808021; 
ram[86]=32'h263128a0; 
ram[87]=32'h8e060000; 
ram[88]=32'h02002821; 
ram[89]=32'h02202021; 
ram[90]=32'h26100004; 
ram[91]=32'h0fc00254; 
ram[92]=32'h00000000; 
ram[93]=32'h1612fff9; 
ram[94]=32'h00000000; 
ram[95]=32'h8fbf001c; 
ram[96]=32'h8fb20018; 
ram[97]=32'h8fb10014; 
ram[98]=32'h8fb00010; 
ram[99]=32'h27bd0020; 
ram[100]=32'h03e00008; 
ram[101]=32'h00000000; 
ram[102]=32'h27bdffc8; 
ram[103]=32'hafb7002c; 
ram[104]=32'hafb60028; 
ram[105]=32'hafb40020; 
ram[106]=32'hafb3001c; 
ram[107]=32'hafb20018; 
ram[108]=32'hafbf0034; 
ram[109]=32'hafbe0030; 
ram[110]=32'hafb50024; 
ram[111]=32'hafb10014; 
ram[112]=32'hafb00010; 
ram[113]=32'h3c179f00; 
ram[114]=32'h0fc0022f; 
ram[115]=32'h00000000; 
ram[116]=32'h3c169f00; 
ram[117]=32'h2413000b; 
ram[118]=32'h2414000c; 
ram[119]=32'h24120001; 
ram[120]=32'h0fc00274; 
ram[121]=32'h00000000; 
ram[122]=32'h10530019; 
ram[123]=32'h00000000; 
ram[124]=32'h1454fffb; 
ram[125]=32'h00000000; 
ram[126]=32'h3c049f00; 
ram[127]=32'h248428e4; 
ram[128]=32'h0fc00254; 
ram[129]=32'h00000000; 
ram[130]=32'h0fc00263; 
ram[131]=32'h00000000; 
ram[132]=32'h3c049f00; 
ram[133]=32'h248428f0; 
ram[134]=32'h00402821; 
ram[135]=32'h00408021; 
ram[136]=32'h0fc00254; 
ram[137]=32'h00000000; 
ram[138]=32'h0fc0023e; 
ram[139]=32'h00000000; 
ram[140]=32'h1452fffd; 
ram[141]=32'h00000000; 
ram[142]=32'h0200f809; 
ram[143]=32'h00000000; 
ram[144]=32'h0fc00274; 
ram[145]=32'h00000000; 
ram[146]=32'h1453ffe9; 
ram[147]=32'h00000000; 
ram[148]=32'h26e428b0; 
ram[149]=32'h0fc00254; 
ram[150]=32'h00000000; 
ram[151]=32'h0fc00263; 
ram[152]=32'h00000000; 
ram[153]=32'h00402821; 
ram[154]=32'h26c428c8; 
ram[155]=32'h00408021; 
ram[156]=32'h0fc00254; 
ram[157]=32'h00000000; 
ram[158]=32'h0fc00263; 
ram[159]=32'h00000000; 
ram[160]=32'h00408821; 
ram[161]=32'h3c029f00; 
ram[162]=32'h244428d8; 
ram[163]=32'h02202821; 
ram[164]=32'h0fc00254; 
ram[165]=32'h00000000; 
ram[166]=32'h1200ffd1; 
ram[167]=32'h00000000; 
ram[168]=32'h0000a821; 
ram[169]=32'h0000f021; 
ram[170]=32'h0fc00274; 
ram[171]=32'h00000000; 
ram[172]=32'h27de0001; 
ram[173]=32'h02b12021; 
ram[174]=32'ha0820000; 
ram[175]=32'h03c0a821; 
ram[176]=32'h17d0fff9; 
ram[177]=32'h00000000; 
ram[178]=32'h0bc00078; 
ram[179]=32'h00000000; 
ram[180]=32'h27bdffe0; 
ram[181]=32'hafb00018; 
ram[182]=32'h3c109f00; 
ram[183]=32'h00002021; 
ram[184]=32'h26052de8; 
ram[185]=32'hafbf001c; 
ram[186]=32'h0fc00394; 
ram[187]=32'h00000000; 
ram[188]=32'h26022de8; 
ram[189]=32'h3c039f00; 
ram[190]=32'h24632be0; 
ram[191]=32'h24440200; 
ram[192]=32'h8c480000; 
ram[193]=32'h8c470004; 
ram[194]=32'h8c460008; 
ram[195]=32'h8c45000c; 
ram[196]=32'h24420010; 
ram[197]=32'hac680000; 
ram[198]=32'hac670004; 
ram[199]=32'hac660008; 
ram[200]=32'hac65000c; 
ram[201]=32'h24630010; 
ram[202]=32'h1444fff5; 
ram[203]=32'h00000000; 
ram[204]=32'h8c440000; 
ram[205]=32'h8fbf001c; 
ram[206]=32'h8c420004; 
ram[207]=32'h8fb00018; 
ram[208]=32'hac620004; 
ram[209]=32'h00001021; 
ram[210]=32'hac640000; 
ram[211]=32'h27bd0020; 
ram[212]=32'h03e00008; 
ram[213]=32'h00000000; 
ram[214]=32'h27bdffc0; 
ram[215]=32'h3c029f00; 
ram[216]=32'h24422be0; 
ram[217]=32'hafbe0038; 
ram[218]=32'hafb70034; 
ram[219]=32'hafb60030; 
ram[220]=32'hafb5002c; 
ram[221]=32'hafb40028; 
ram[222]=32'hafb30024; 
ram[223]=32'hafb20020; 
ram[224]=32'hafb1001c; 
ram[225]=32'hafb00018; 
ram[226]=32'hafbf003c; 
ram[227]=32'h8c430030; 
ram[228]=32'h9045000e; 
ram[229]=32'h2463fffe; 
ram[230]=32'h00a30018; 
ram[231]=32'h90460012; 
ram[232]=32'h8c450028; 
ram[233]=32'h94430010; 
ram[234]=32'h70c50000; 
ram[235]=32'h944a000c; 
ram[236]=32'h00002812; 
ram[237]=32'h3c119f00; 
ram[238]=32'h00a31021; 
ram[239]=32'h71429802; 
ram[240]=32'h26302de8; 
ram[241]=32'h3c099f00; 
ram[242]=32'h0080b021; 
ram[243]=32'h0000a821; 
ram[244]=32'h261e0200; 
ram[245]=32'h3c179f00; 
ram[246]=32'h25322960; 
ram[247]=32'h2414000b; 
ram[248]=32'h2a620000; 
ram[249]=32'h266401ff; 
ram[250]=32'h0262200a; 
ram[251]=32'h00042243; 
ram[252]=32'h02002821; 
ram[253]=32'h0fc00394; 
ram[254]=32'h00000000; 
ram[255]=32'h92222de8; 
ram[256]=32'h10400036; 
ram[257]=32'h00000000; 
ram[258]=32'h3c039f00; 
ram[259]=32'h3c079f00; 
ram[260]=32'h24682e08; 
ram[261]=32'h24e72de8; 
ram[262]=32'h2404000a; 
ram[263]=32'h240b00e5; 
ram[264]=32'h90e3000b; 
ram[265]=32'h30630008; 
ram[266]=32'h10600003; 
ram[267]=32'h00000000; 
ram[268]=32'h104b0023; 
ram[269]=32'h00000000; 
ram[270]=32'h8ee32950; 
ram[271]=32'h8ce5001c; 
ram[272]=32'h00031140; 
ram[273]=32'h8cf90000; 
ram[274]=32'h8cf80004; 
ram[275]=32'h8cef0008; 
ram[276]=32'h8cee000c; 
ram[277]=32'h8ced0010; 
ram[278]=32'h8cec0014; 
ram[279]=32'h8ce60018; 
ram[280]=32'h00521021; 
ram[281]=32'h24630001; 
ram[282]=32'hac45001c; 
ram[283]=32'hac590000; 
ram[284]=32'hac580004; 
ram[285]=32'hac4f0008; 
ram[286]=32'hac4e000c; 
ram[287]=32'hac4d0010; 
ram[288]=32'hac4c0014; 
ram[289]=32'hac460018; 
ram[290]=32'haee32950; 
ram[291]=32'h00001021; 
ram[292]=32'h02d52821; 
ram[293]=32'h00e21821; 
ram[294]=32'h90660000; 
ram[295]=32'h00a21821; 
ram[296]=32'h24420001; 
ram[297]=32'ha0660000; 
ram[298]=32'h1454fffa; 
ram[299]=32'h00000000; 
ram[300]=32'h26a2000b; 
ram[301]=32'h02c21021; 
ram[302]=32'h26b5000c; 
ram[303]=32'ha0440000; 
ram[304]=32'h111e0016; 
ram[305]=32'h00000000; 
ram[306]=32'h01003821; 
ram[307]=32'h25080020; 
ram[308]=32'h9102ffe0; 
ram[309]=32'h1440ffd2; 
ram[310]=32'h00000000; 
ram[311]=32'h02d5a821; 
ram[312]=32'ha2a00000; 
ram[313]=32'h8fbf003c; 
ram[314]=32'h8fbe0038; 
ram[315]=32'h8fb70034; 
ram[316]=32'h8fb60030; 
ram[317]=32'h8fb5002c; 
ram[318]=32'h8fb40028; 
ram[319]=32'h8fb30024; 
ram[320]=32'h8fb20020; 
ram[321]=32'h8fb1001c; 
ram[322]=32'h8fb00018; 
ram[323]=32'h00001021; 
ram[324]=32'h27bd0040; 
ram[325]=32'h03e00008; 
ram[326]=32'h00000000; 
ram[327]=32'h26730200; 
ram[328]=32'h0bc000f8; 
ram[329]=32'h00000000; 
ram[330]=32'h3c029f00; 
ram[331]=32'h8c462950; 
ram[332]=32'h10c00034; 
ram[333]=32'h00000000; 
ram[334]=32'h3c039f00; 
ram[335]=32'h24632960; 
ram[336]=32'h00001021; 
ram[337]=32'h0bc00157; 
ram[338]=32'h00000000; 
ram[339]=32'h24420001; 
ram[340]=32'h24630020; 
ram[341]=32'h1046002b; 
ram[342]=32'h00000000; 
ram[343]=32'h9065000b; 
ram[344]=32'h30a50018; 
ram[345]=32'h14a0fff9; 
ram[346]=32'h00000000; 
ram[347]=32'h00003021; 
ram[348]=32'h00004021; 
ram[349]=32'h24090020; 
ram[350]=32'h240b007e; 
ram[351]=32'h240d0031; 
ram[352]=32'h240a0008; 
ram[353]=32'h90650000; 
ram[354]=32'h10a90019; 
ram[355]=32'h00000000; 
ram[356]=32'h10ab0010; 
ram[357]=32'h00000000; 
ram[358]=32'h90870000; 
ram[359]=32'h10a70006; 
ram[360]=32'h00000000; 
ram[361]=32'h24a50020; 
ram[362]=32'h10a70003; 
ram[363]=32'h00000000; 
ram[364]=32'h15000015; 
ram[365]=32'h00000000; 
ram[366]=32'h24c60001; 
ram[367]=32'h24630001; 
ram[368]=32'h24840001; 
ram[369]=32'h14caffef; 
ram[370]=32'h00000000; 
ram[371]=32'h03e00008; 
ram[372]=32'h00000000; 
ram[373]=32'h90670001; 
ram[374]=32'h14edffef; 
ram[375]=32'h00000000; 
ram[376]=32'h90870000; 
ram[377]=32'h24080001; 
ram[378]=32'h0bc00167; 
ram[379]=32'h00000000; 
ram[380]=32'h90870000; 
ram[381]=32'h240c0001; 
ram[382]=32'h0187400a; 
ram[383]=32'h0bc00167; 
ram[384]=32'h00000000; 
ram[385]=32'h2402ffff; 
ram[386]=32'h03e00008; 
ram[387]=32'h00000000; 
ram[388]=32'h27bdffe0; 
ram[389]=32'hafbf001c; 
ram[390]=32'h0fc0014a; 
ram[391]=32'h00000000; 
ram[392]=32'h0440000a; 
ram[393]=32'h00000000; 
ram[394]=32'h3c039f00; 
ram[395]=32'h00021140; 
ram[396]=32'h24632960; 
ram[397]=32'h00621021; 
ram[398]=32'h8c42001c; 
ram[399]=32'h8fbf001c; 
ram[400]=32'h27bd0020; 
ram[401]=32'h03e00008; 
ram[402]=32'h00000000; 
ram[403]=32'h2402ffff; 
ram[404]=32'h0bc0018f; 
ram[405]=32'h00000000; 
ram[406]=32'h27bdffc8; 
ram[407]=32'h00a07021; 
ram[408]=32'hafb60030; 
ram[409]=32'hafb5002c; 
ram[410]=32'hafbf0034; 
ram[411]=32'hafb40028; 
ram[412]=32'hafb30024; 
ram[413]=32'hafb20020; 
ram[414]=32'hafb1001c; 
ram[415]=32'hafb00018; 
ram[416]=32'h00c0b021; 
ram[417]=32'h00e0a821; 
ram[418]=32'h0fc0014a; 
ram[419]=32'h00000000; 
ram[420]=32'h0440004d; 
ram[421]=32'h00000000; 
ram[422]=32'h3c039f00; 
ram[423]=32'h00021140; 
ram[424]=32'h24632960; 
ram[425]=32'h00431821; 
ram[426]=32'h3c029f00; 
ram[427]=32'h24422be0; 
ram[428]=32'h94650014; 
ram[429]=32'h94470010; 
ram[430]=32'h9464001a; 
ram[431]=32'h90460012; 
ram[432]=32'h8c430028; 
ram[433]=32'h00052c00; 
ram[434]=32'h00e00013; 
ram[435]=32'h00a42821; 
ram[436]=32'h70c30000; 
ram[437]=32'h9044000e; 
ram[438]=32'h24a5fffc; 
ram[439]=32'h70a40000; 
ram[440]=32'h9443000c; 
ram[441]=32'h00001012; 
ram[442]=32'h70622002; 
ram[443]=32'h008e1021; 
ram[444]=32'h1ac0001f; 
ram[445]=32'h00000000; 
ram[446]=32'h244301ff; 
ram[447]=32'h28440000; 
ram[448]=32'h0064100b; 
ram[449]=32'h3c119f00; 
ram[450]=32'h00029a43; 
ram[451]=32'h26252de8; 
ram[452]=32'h02602021; 
ram[453]=32'h00a09021; 
ram[454]=32'h0240a021; 
ram[455]=32'h0fc00394; 
ram[456]=32'h00000000; 
ram[457]=32'h00002021; 
ram[458]=32'h92232de8; 
ram[459]=32'h02a41021; 
ram[460]=32'h24900001; 
ram[461]=32'h24850200; 
ram[462]=32'ha0430000; 
ram[463]=32'h02442023; 
ram[464]=32'h0bc001d6; 
ram[465]=32'h00000000; 
ram[466]=32'h9102ffff; 
ram[467]=32'ha062ffff; 
ram[468]=32'h12050013; 
ram[469]=32'h00000000; 
ram[470]=32'h0216102a; 
ram[471]=32'h26100001; 
ram[472]=32'h00904021; 
ram[473]=32'h02b01821; 
ram[474]=32'h1440fff7; 
ram[475]=32'h00000000; 
ram[476]=32'h00001021; 
ram[477]=32'h8fbf0034; 
ram[478]=32'h8fb60030; 
ram[479]=32'h8fb5002c; 
ram[480]=32'h8fb40028; 
ram[481]=32'h8fb30024; 
ram[482]=32'h8fb20020; 
ram[483]=32'h8fb1001c; 
ram[484]=32'h8fb00018; 
ram[485]=32'h27bd0038; 
ram[486]=32'h03e00008; 
ram[487]=32'h00000000; 
ram[488]=32'h0216102a; 
ram[489]=32'h1040fff2; 
ram[490]=32'h00000000; 
ram[491]=32'h02602021; 
ram[492]=32'h02802821; 
ram[493]=32'h0fc00394; 
ram[494]=32'h00000000; 
ram[495]=32'h02002021; 
ram[496]=32'h0bc001ca; 
ram[497]=32'h00000000; 
ram[498]=32'h2402ffff; 
ram[499]=32'h0bc001dd; 
ram[500]=32'h00000000; 
ram[501]=32'h00000000; 
ram[502]=32'h00000000; 
ram[503]=32'h00000000; 
ram[504]=32'h3c02b801; 
ram[505]=32'ha04012c0; 
ram[506]=32'h03e00008; 
ram[507]=32'h00000000; 
ram[508]=32'h00063600; 
ram[509]=32'h2c82003d; 
ram[510]=32'h00063603; 
ram[511]=32'h1040000c; 
ram[512]=32'h00000000; 
ram[513]=32'h2ca20051; 
ram[514]=32'h10400009; 
ram[515]=32'h00000000; 
ram[516]=32'h00041100; 
ram[517]=32'h00042180; 
ram[518]=32'h00442021; 
ram[519]=32'h00852821; 
ram[520]=32'h3c02b801; 
ram[521]=32'h30c600ff; 
ram[522]=32'h00a22821; 
ram[523]=32'ha0a60000; 
ram[524]=32'h03e00008; 
ram[525]=32'h00000000; 
ram[526]=32'h00041900; 
ram[527]=32'h80c20000; 
ram[528]=32'h00042180; 
ram[529]=32'h00642021; 
ram[530]=32'h00852821; 
ram[531]=32'h1040000b; 
ram[532]=32'h00000000; 
ram[533]=32'h3c04b801; 
ram[534]=32'h00862023; 
ram[535]=32'h00852021; 
ram[536]=32'h00c41821; 
ram[537]=32'h304200ff; 
ram[538]=32'ha0620000; 
ram[539]=32'h24c60001; 
ram[540]=32'h80c20000; 
ram[541]=32'h1440fffa; 
ram[542]=32'h00000000; 
ram[543]=32'h03e00008; 
ram[544]=32'h00000000; 
ram[545]=32'h00000000; 
ram[546]=32'h00000000; 
ram[547]=32'h00000000; 
ram[548]=32'h00042600; 
ram[549]=32'h00042603; 
ram[550]=32'h3c02b800; 
ram[551]=32'h904303fd; 
ram[552]=32'h30630020; 
ram[553]=32'h1060fffc; 
ram[554]=32'h00000000; 
ram[555]=32'h308300ff; 
ram[556]=32'ha04303f8; 
ram[557]=32'h03e00008; 
ram[558]=32'h00000000; 
ram[559]=32'h3c02b800; 
ram[560]=32'h2403ff80; 
ram[561]=32'ha04003f9; 
ram[562]=32'ha04303fb; 
ram[563]=32'h2403001b; 
ram[564]=32'ha04303f8; 
ram[565]=32'h24030003; 
ram[566]=32'ha04003f9; 
ram[567]=32'ha04303fb; 
ram[568]=32'h2403ffc7; 
ram[569]=32'ha04303fa; 
ram[570]=32'h2403000b; 
ram[571]=32'ha04303fc; 
ram[572]=32'h03e00008; 
ram[573]=32'h00000000; 
ram[574]=32'h3c02b800; 
ram[575]=32'h904203fd; 
ram[576]=32'h00021142; 
ram[577]=32'h30420001; 
ram[578]=32'h03e00008; 
ram[579]=32'h00000000; 
ram[580]=32'h80860000; 
ram[581]=32'h3c02b800; 
ram[582]=32'h10c0000b; 
ram[583]=32'h00000000; 
ram[584]=32'h904303fd; 
ram[585]=32'h30630020; 
ram[586]=32'h1060fffd; 
ram[587]=32'h00000000; 
ram[588]=32'h30c600ff; 
ram[589]=32'ha04603f8; 
ram[590]=32'h24840001; 
ram[591]=32'h80860000; 
ram[592]=32'h14c0fff7; 
ram[593]=32'h00000000; 
ram[594]=32'h03e00008; 
ram[595]=32'h00000000; 
ram[596]=32'h27bdffe0; 
ram[597]=32'hafa60028; 
ram[598]=32'h3c069f00; 
ram[599]=32'hafa50024; 
ram[600]=32'h24c60890; 
ram[601]=32'h27a50024; 
ram[602]=32'hafbf001c; 
ram[603]=32'hafa7002c; 
ram[604]=32'hafa40020; 
ram[605]=32'h0fc00979; 
ram[606]=32'h00000000; 
ram[607]=32'h8fbf001c; 
ram[608]=32'h27bd0020; 
ram[609]=32'h03e00008; 
ram[610]=32'h00000000; 
ram[611]=32'h00003021; 
ram[612]=32'h00001021; 
ram[613]=32'h3c03b800; 
ram[614]=32'h24070020; 
ram[615]=32'h906403fd; 
ram[616]=32'h30840001; 
ram[617]=32'h1080fffd; 
ram[618]=32'h00000000; 
ram[619]=32'h906403f8; 
ram[620]=32'h308400ff; 
ram[621]=32'h00c42004; 
ram[622]=32'h24c60008; 
ram[623]=32'h00441025; 
ram[624]=32'h14c7fff6; 
ram[625]=32'h00000000; 
ram[626]=32'h03e00008; 
ram[627]=32'h00000000; 
ram[628]=32'h3c02b800; 
ram[629]=32'h904303fd; 
ram[630]=32'h30630001; 
ram[631]=32'h1060fffc; 
ram[632]=32'h00000000; 
ram[633]=32'h904203f8; 
ram[634]=32'h304200ff; 
ram[635]=32'h03e00008; 
ram[636]=32'h00000000; 
ram[637]=32'h18a0000c; 
ram[638]=32'h00000000; 
ram[639]=32'h00853021; 
ram[640]=32'h3c02b800; 
ram[641]=32'h904303fd; 
ram[642]=32'h30630001; 
ram[643]=32'h1060fffd; 
ram[644]=32'h00000000; 
ram[645]=32'h904303f8; 
ram[646]=32'h24840001; 
ram[647]=32'ha083ffff; 
ram[648]=32'h1486fff8; 
ram[649]=32'h00000000; 
ram[650]=32'h03e00008; 
ram[651]=32'h00000000; 
ram[652]=32'h3c02b800; 
ram[653]=32'h2403ffff; 
ram[654]=32'hac440404; 
ram[655]=32'hac430400; 
ram[656]=32'h03e00008; 
ram[657]=32'h00000000; 
ram[658]=32'h3c02b800; 
ram[659]=32'h8c430400; 
ram[660]=32'h24050001; 
ram[661]=32'h00852004; 
ram[662]=32'h00831825; 
ram[663]=32'hac430400; 
ram[664]=32'h03e00008; 
ram[665]=32'h00000000; 
ram[666]=32'h3c02b800; 
ram[667]=32'h24050001; 
ram[668]=32'h8c430400; 
ram[669]=32'h00852004; 
ram[670]=32'h00042827; 
ram[671]=32'h00a31824; 
ram[672]=32'hac430400; 
ram[673]=32'h03e00008; 
ram[674]=32'h00000000; 
ram[675]=32'h3c02b800; 
ram[676]=32'h8c430400; 
ram[677]=32'h24020001; 
ram[678]=32'h00821004; 
ram[679]=32'h00431024; 
ram[680]=32'h03e00008; 
ram[681]=32'h00000000; 
ram[682]=32'h00000000; 
ram[683]=32'h00000000; 
ram[684]=32'h308400ff; 
ram[685]=32'h0bc005e9; 
ram[686]=32'h00000000; 
ram[687]=32'h240400ff; 
ram[688]=32'h0bc005e9; 
ram[689]=32'h00000000; 
ram[690]=32'h00002021; 
ram[691]=32'h0bc005f5; 
ram[692]=32'h00000000; 
ram[693]=32'h27bdffe0; 
ram[694]=32'hafbf001c; 
ram[695]=32'h0fc005fd; 
ram[696]=32'h00000000; 
ram[697]=32'h8fbf001c; 
ram[698]=32'h240400ff; 
ram[699]=32'h27bd0020; 
ram[700]=32'h0bc005e9; 
ram[701]=32'h00000000; 
ram[702]=32'h27bdffd8; 
ram[703]=32'h3084003f; 
ram[704]=32'h34840040; 
ram[705]=32'hafb0001c; 
ram[706]=32'h00a08021; 
ram[707]=32'hafbf0024; 
ram[708]=32'hafb10020; 
ram[709]=32'h30d100ff; 
ram[710]=32'h0fc005e9; 
ram[711]=32'h00000000; 
ram[712]=32'h00102602; 
ram[713]=32'h0fc005e9; 
ram[714]=32'h00000000; 
ram[715]=32'h00102402; 
ram[716]=32'h308400ff; 
ram[717]=32'h0fc005e9; 
ram[718]=32'h00000000; 
ram[719]=32'h00102202; 
ram[720]=32'h308400ff; 
ram[721]=32'h0fc005e9; 
ram[722]=32'h00000000; 
ram[723]=32'h320400ff; 
ram[724]=32'h0fc005e9; 
ram[725]=32'h00000000; 
ram[726]=32'h02202021; 
ram[727]=32'h0fc005e9; 
ram[728]=32'h00000000; 
ram[729]=32'h240400ff; 
ram[730]=32'h241000fe; 
ram[731]=32'h0fc005e9; 
ram[732]=32'h00000000; 
ram[733]=32'h241100ff; 
ram[734]=32'h0bc002e6; 
ram[735]=32'h00000000; 
ram[736]=32'h2610ffff; 
ram[737]=32'h321000ff; 
ram[738]=32'h0fc005e9; 
ram[739]=32'h00000000; 
ram[740]=32'h12000004; 
ram[741]=32'h00000000; 
ram[742]=32'h240400ff; 
ram[743]=32'h1051fff8; 
ram[744]=32'h00000000; 
ram[745]=32'h8fbf0024; 
ram[746]=32'h8fb10020; 
ram[747]=32'h8fb0001c; 
ram[748]=32'h27bd0028; 
ram[749]=32'h03e00008; 
ram[750]=32'h00000000; 
ram[751]=32'h27bdffd0; 
ram[752]=32'hafbf002c; 
ram[753]=32'hafb10024; 
ram[754]=32'hafb20028; 
ram[755]=32'hafb00020; 
ram[756]=32'h24110010; 
ram[757]=32'h0fc005fd; 
ram[758]=32'h00000000; 
ram[759]=32'h240400ff; 
ram[760]=32'h0fc005e9; 
ram[761]=32'h00000000; 
ram[762]=32'h2631ffff; 
ram[763]=32'h240400ff; 
ram[764]=32'h323100ff; 
ram[765]=32'h0fc005e9; 
ram[766]=32'h00000000; 
ram[767]=32'h1620fffa; 
ram[768]=32'h00000000; 
ram[769]=32'h00002021; 
ram[770]=32'h0fc005f5; 
ram[771]=32'h00000000; 
ram[772]=32'h00002021; 
ram[773]=32'h00002821; 
ram[774]=32'h24060095; 
ram[775]=32'h241000fe; 
ram[776]=32'h0fc002be; 
ram[777]=32'h00000000; 
ram[778]=32'h24120001; 
ram[779]=32'h0bc00313; 
ram[780]=32'h00000000; 
ram[781]=32'h2610ffff; 
ram[782]=32'h321000ff; 
ram[783]=32'h0fc002be; 
ram[784]=32'h00000000; 
ram[785]=32'h12000013; 
ram[786]=32'h00000000; 
ram[787]=32'h00002021; 
ram[788]=32'h00002821; 
ram[789]=32'h24060095; 
ram[790]=32'h1452fff6; 
ram[791]=32'h00000000; 
ram[792]=32'h0fc005fd; 
ram[793]=32'h00000000; 
ram[794]=32'h240400ff; 
ram[795]=32'h0fc005e9; 
ram[796]=32'h00000000; 
ram[797]=32'h8fbf002c; 
ram[798]=32'h02201021; 
ram[799]=32'h8fb20028; 
ram[800]=32'h8fb10024; 
ram[801]=32'h8fb00020; 
ram[802]=32'h27bd0030; 
ram[803]=32'h03e00008; 
ram[804]=32'h00000000; 
ram[805]=32'hafa20018; 
ram[806]=32'h0fc005fd; 
ram[807]=32'h00000000; 
ram[808]=32'h8fa20018; 
ram[809]=32'h240400ff; 
ram[810]=32'h00408821; 
ram[811]=32'h0fc005e9; 
ram[812]=32'h00000000; 
ram[813]=32'h8fbf002c; 
ram[814]=32'h02201021; 
ram[815]=32'h8fb20028; 
ram[816]=32'h8fb10024; 
ram[817]=32'h8fb00020; 
ram[818]=32'h27bd0030; 
ram[819]=32'h03e00008; 
ram[820]=32'h00000000; 
ram[821]=32'h27bdffd0; 
ram[822]=32'h00002021; 
ram[823]=32'hafbf002c; 
ram[824]=32'hafb30028; 
ram[825]=32'hafb20024; 
ram[826]=32'hafb10020; 
ram[827]=32'hafb0001c; 
ram[828]=32'h0fc005f5; 
ram[829]=32'h00000000; 
ram[830]=32'h24040008; 
ram[831]=32'h240501aa; 
ram[832]=32'h24060087; 
ram[833]=32'h0fc002be; 
ram[834]=32'h00000000; 
ram[835]=32'h24030005; 
ram[836]=32'h10430041; 
ram[837]=32'h00000000; 
ram[838]=32'h240400ff; 
ram[839]=32'h0fc005e9; 
ram[840]=32'h00000000; 
ram[841]=32'h240400ff; 
ram[842]=32'h0fc005e9; 
ram[843]=32'h00000000; 
ram[844]=32'h240400ff; 
ram[845]=32'h0fc005e9; 
ram[846]=32'h00000000; 
ram[847]=32'h240400ff; 
ram[848]=32'h00008021; 
ram[849]=32'h0fc005e9; 
ram[850]=32'h00000000; 
ram[851]=32'h24130001; 
ram[852]=32'h0bc00359; 
ram[853]=32'h00000000; 
ram[854]=32'h1053001b; 
ram[855]=32'h00000000; 
ram[856]=32'h00608021; 
ram[857]=32'h24040037; 
ram[858]=32'h00002821; 
ram[859]=32'h240600ff; 
ram[860]=32'h0fc002be; 
ram[861]=32'h00000000; 
ram[862]=32'h26030001; 
ram[863]=32'h306300ff; 
ram[864]=32'h241100ff; 
ram[865]=32'h00409021; 
ram[866]=32'h1471fff3; 
ram[867]=32'h00000000; 
ram[868]=32'h0fc005fd; 
ram[869]=32'h00000000; 
ram[870]=32'h240400ff; 
ram[871]=32'h0fc005e9; 
ram[872]=32'h00000000; 
ram[873]=32'h02401021; 
ram[874]=32'h8fbf002c; 
ram[875]=32'h8fb30028; 
ram[876]=32'h8fb20024; 
ram[877]=32'h8fb10020; 
ram[878]=32'h8fb0001c; 
ram[879]=32'h27bd0030; 
ram[880]=32'h03e00008; 
ram[881]=32'h00000000; 
ram[882]=32'h24040029; 
ram[883]=32'h3c054000; 
ram[884]=32'h240600ff; 
ram[885]=32'h26100002; 
ram[886]=32'h0fc002be; 
ram[887]=32'h00000000; 
ram[888]=32'h321000ff; 
ram[889]=32'h00409021; 
ram[890]=32'h1211ffe9; 
ram[891]=32'h00000000; 
ram[892]=32'h1440ffdc; 
ram[893]=32'h00000000; 
ram[894]=32'h0fc005fd; 
ram[895]=32'h00000000; 
ram[896]=32'h240400ff; 
ram[897]=32'h0fc005e9; 
ram[898]=32'h00000000; 
ram[899]=32'h00001021; 
ram[900]=32'h0bc0036a; 
ram[901]=32'h00000000; 
ram[902]=32'h0fc005fd; 
ram[903]=32'h00000000; 
ram[904]=32'h240400ff; 
ram[905]=32'h0fc005e9; 
ram[906]=32'h00000000; 
ram[907]=32'h8fbf002c; 
ram[908]=32'h8fb30028; 
ram[909]=32'h8fb20024; 
ram[910]=32'h8fb10020; 
ram[911]=32'h8fb0001c; 
ram[912]=32'h24020005; 
ram[913]=32'h27bd0030; 
ram[914]=32'h03e00008; 
ram[915]=32'h00000000; 
ram[916]=32'h27bdffc8; 
ram[917]=32'hafb00024; 
ram[918]=32'h00808021; 
ram[919]=32'h00002021; 
ram[920]=32'hafbf0034; 
ram[921]=32'hafb10028; 
ram[922]=32'hafb30030; 
ram[923]=32'h00a08821; 
ram[924]=32'hafb2002c; 
ram[925]=32'h0fc005f5; 
ram[926]=32'h00000000; 
ram[927]=32'h24040011; 
ram[928]=32'h00102a40; 
ram[929]=32'h24060055; 
ram[930]=32'h0fc002be; 
ram[931]=32'h00000000; 
ram[932]=32'h14400032; 
ram[933]=32'h00000000; 
ram[934]=32'h240400ff; 
ram[935]=32'h0fc005e9; 
ram[936]=32'h00000000; 
ram[937]=32'h00409021; 
ram[938]=32'h24107530; 
ram[939]=32'h241300fe; 
ram[940]=32'h0bc003b5; 
ram[941]=32'h00000000; 
ram[942]=32'h2610ffff; 
ram[943]=32'h0fc005e9; 
ram[944]=32'h00000000; 
ram[945]=32'h3210ffff; 
ram[946]=32'h00409021; 
ram[947]=32'h12000034; 
ram[948]=32'h00000000; 
ram[949]=32'h240400ff; 
ram[950]=32'h1653fff7; 
ram[951]=32'h00000000; 
ram[952]=32'h00008021; 
ram[953]=32'h24120200; 
ram[954]=32'h240400ff; 
ram[955]=32'h0fc005e9; 
ram[956]=32'h00000000; 
ram[957]=32'h02301821; 
ram[958]=32'h26100001; 
ram[959]=32'ha0620000; 
ram[960]=32'h1612fff9; 
ram[961]=32'h00000000; 
ram[962]=32'h240400ff; 
ram[963]=32'h0fc005e9; 
ram[964]=32'h00000000; 
ram[965]=32'h240400ff; 
ram[966]=32'h0fc005e9; 
ram[967]=32'h00000000; 
ram[968]=32'h0fc005fd; 
ram[969]=32'h00000000; 
ram[970]=32'h240400ff; 
ram[971]=32'h0fc005e9; 
ram[972]=32'h00000000; 
ram[973]=32'h8fbf0034; 
ram[974]=32'h00009021; 
ram[975]=32'h02401021; 
ram[976]=32'h8fb30030; 
ram[977]=32'h8fb2002c; 
ram[978]=32'h8fb10028; 
ram[979]=32'h8fb00024; 
ram[980]=32'h27bd0038; 
ram[981]=32'h03e00008; 
ram[982]=32'h00000000; 
ram[983]=32'hafa20018; 
ram[984]=32'h0fc005fd; 
ram[985]=32'h00000000; 
ram[986]=32'h8fa20018; 
ram[987]=32'h240400ff; 
ram[988]=32'h00409021; 
ram[989]=32'h0fc005e9; 
ram[990]=32'h00000000; 
ram[991]=32'h8fbf0034; 
ram[992]=32'h02401021; 
ram[993]=32'h8fb30030; 
ram[994]=32'h8fb2002c; 
ram[995]=32'h8fb10028; 
ram[996]=32'h8fb00024; 
ram[997]=32'h27bd0038; 
ram[998]=32'h03e00008; 
ram[999]=32'h00000000; 
ram[1000]=32'h0fc005fd; 
ram[1001]=32'h00000000; 
ram[1002]=32'h240400ff; 
ram[1003]=32'h0fc005e9; 
ram[1004]=32'h00000000; 
ram[1005]=32'h8fbf0034; 
ram[1006]=32'h02401021; 
ram[1007]=32'h8fb30030; 
ram[1008]=32'h8fb2002c; 
ram[1009]=32'h8fb10028; 
ram[1010]=32'h8fb00024; 
ram[1011]=32'h27bd0038; 
ram[1012]=32'h03e00008; 
ram[1013]=32'h00000000; 
ram[1014]=32'h27bdffc8; 
ram[1015]=32'hafb10024; 
ram[1016]=32'h00808821; 
ram[1017]=32'h00002021; 
ram[1018]=32'hafbf0034; 
ram[1019]=32'hafb40030; 
ram[1020]=32'hafb00020; 
ram[1021]=32'h30b400ff; 
ram[1022]=32'h00c08021; 
ram[1023]=32'hafb3002c; 
ram[1024]=32'hafb20028; 
ram[1025]=32'h0fc005f5; 
ram[1026]=32'h00000000; 
ram[1027]=32'h24040012; 
ram[1028]=32'h00112a40; 
ram[1029]=32'h240600ff; 
ram[1030]=32'h0fc002be; 
ram[1031]=32'h00000000; 
ram[1032]=32'h1440003f; 
ram[1033]=32'h00000000; 
ram[1034]=32'h241300fe; 
ram[1035]=32'h240400ff; 
ram[1036]=32'h0fc005e9; 
ram[1037]=32'h00000000; 
ram[1038]=32'h00408821; 
ram[1039]=32'h24127530; 
ram[1040]=32'h0bc0041b; 
ram[1041]=32'h00000000; 
ram[1042]=32'h16200026; 
ram[1043]=32'h00000000; 
ram[1044]=32'h2652ffff; 
ram[1045]=32'h0fc005e9; 
ram[1046]=32'h00000000; 
ram[1047]=32'h3252ffff; 
ram[1048]=32'h00408821; 
ram[1049]=32'h1240001f; 
ram[1050]=32'h00000000; 
ram[1051]=32'h322200f0; 
ram[1052]=32'h240400ff; 
ram[1053]=32'h1040fff4; 
ram[1054]=32'h00000000; 
ram[1055]=32'h1633fff4; 
ram[1056]=32'h00000000; 
ram[1057]=32'h26110200; 
ram[1058]=32'h240400ff; 
ram[1059]=32'h0fc005e9; 
ram[1060]=32'h00000000; 
ram[1061]=32'h26100001; 
ram[1062]=32'ha202ffff; 
ram[1063]=32'h1611fffa; 
ram[1064]=32'h00000000; 
ram[1065]=32'h240400ff; 
ram[1066]=32'h2694ffff; 
ram[1067]=32'h0fc005e9; 
ram[1068]=32'h00000000; 
ram[1069]=32'h329400ff; 
ram[1070]=32'h240400ff; 
ram[1071]=32'h0fc005e9; 
ram[1072]=32'h00000000; 
ram[1073]=32'h1680ffd9; 
ram[1074]=32'h00000000; 
ram[1075]=32'h2404000c; 
ram[1076]=32'h00002821; 
ram[1077]=32'h240600ff; 
ram[1078]=32'h00008821; 
ram[1079]=32'h0fc002be; 
ram[1080]=32'h00000000; 
ram[1081]=32'h0fc005fd; 
ram[1082]=32'h00000000; 
ram[1083]=32'h240400ff; 
ram[1084]=32'h0fc005e9; 
ram[1085]=32'h00000000; 
ram[1086]=32'h8fbf0034; 
ram[1087]=32'h02201021; 
ram[1088]=32'h8fb40030; 
ram[1089]=32'h8fb3002c; 
ram[1090]=32'h8fb20028; 
ram[1091]=32'h8fb10024; 
ram[1092]=32'h8fb00020; 
ram[1093]=32'h27bd0038; 
ram[1094]=32'h03e00008; 
ram[1095]=32'h00000000; 
ram[1096]=32'hafa20018; 
ram[1097]=32'h0fc005fd; 
ram[1098]=32'h00000000; 
ram[1099]=32'h8fa20018; 
ram[1100]=32'h240400ff; 
ram[1101]=32'h00408821; 
ram[1102]=32'h0fc005e9; 
ram[1103]=32'h00000000; 
ram[1104]=32'h8fbf0034; 
ram[1105]=32'h02201021; 
ram[1106]=32'h8fb40030; 
ram[1107]=32'h8fb3002c; 
ram[1108]=32'h8fb20028; 
ram[1109]=32'h8fb10024; 
ram[1110]=32'h8fb00020; 
ram[1111]=32'h27bd0038; 
ram[1112]=32'h03e00008; 
ram[1113]=32'h00000000; 
ram[1114]=32'h27bdffc8; 
ram[1115]=32'hafb30030; 
ram[1116]=32'h00049a40; 
ram[1117]=32'h00002021; 
ram[1118]=32'hafb2002c; 
ram[1119]=32'hafb10028; 
ram[1120]=32'hafb00024; 
ram[1121]=32'hafbf0034; 
ram[1122]=32'h00a08821; 
ram[1123]=32'h00008021; 
ram[1124]=32'h0fc005f5; 
ram[1125]=32'h00000000; 
ram[1126]=32'h24120200; 
ram[1127]=32'h0bc0046b; 
ram[1128]=32'h00000000; 
ram[1129]=32'h1040001c; 
ram[1130]=32'h00000000; 
ram[1131]=32'h26100001; 
ram[1132]=32'h24040018; 
ram[1133]=32'h02602821; 
ram[1134]=32'h240600ff; 
ram[1135]=32'h3210ffff; 
ram[1136]=32'h0fc002be; 
ram[1137]=32'h00000000; 
ram[1138]=32'h2e0300ff; 
ram[1139]=32'h1460fff5; 
ram[1140]=32'h00000000; 
ram[1141]=32'hafa20018; 
ram[1142]=32'h0fc005fd; 
ram[1143]=32'h00000000; 
ram[1144]=32'h8fa20018; 
ram[1145]=32'h240400ff; 
ram[1146]=32'h00408021; 
ram[1147]=32'h0fc005e9; 
ram[1148]=32'h00000000; 
ram[1149]=32'h8fbf0034; 
ram[1150]=32'h02001021; 
ram[1151]=32'h8fb30030; 
ram[1152]=32'h8fb2002c; 
ram[1153]=32'h8fb10028; 
ram[1154]=32'h8fb00024; 
ram[1155]=32'h27bd0038; 
ram[1156]=32'h03e00008; 
ram[1157]=32'h00000000; 
ram[1158]=32'h24100005; 
ram[1159]=32'h2610ffff; 
ram[1160]=32'h240400ff; 
ram[1161]=32'h3210ffff; 
ram[1162]=32'h0fc005e9; 
ram[1163]=32'h00000000; 
ram[1164]=32'h1600fffa; 
ram[1165]=32'h00000000; 
ram[1166]=32'h240400fe; 
ram[1167]=32'h0fc005e9; 
ram[1168]=32'h00000000; 
ram[1169]=32'h02301021; 
ram[1170]=32'h90440000; 
ram[1171]=32'h26100001; 
ram[1172]=32'h0fc005e9; 
ram[1173]=32'h00000000; 
ram[1174]=32'h1612fffa; 
ram[1175]=32'h00000000; 
ram[1176]=32'h240400ff; 
ram[1177]=32'h0fc005e9; 
ram[1178]=32'h00000000; 
ram[1179]=32'h240400ff; 
ram[1180]=32'h0fc005e9; 
ram[1181]=32'h00000000; 
ram[1182]=32'h240400ff; 
ram[1183]=32'h0fc005e9; 
ram[1184]=32'h00000000; 
ram[1185]=32'h3042001f; 
ram[1186]=32'h24030005; 
ram[1187]=32'h10430004; 
ram[1188]=32'h00000000; 
ram[1189]=32'h24100001; 
ram[1190]=32'h0bc0046b; 
ram[1191]=32'h00000000; 
ram[1192]=32'h240400ff; 
ram[1193]=32'h0fc005e9; 
ram[1194]=32'h00000000; 
ram[1195]=32'h00408021; 
ram[1196]=32'h3411ea60; 
ram[1197]=32'h241200ff; 
ram[1198]=32'h0bc004b7; 
ram[1199]=32'h00000000; 
ram[1200]=32'h2631ffff; 
ram[1201]=32'h0fc005e9; 
ram[1202]=32'h00000000; 
ram[1203]=32'h3231ffff; 
ram[1204]=32'h00408021; 
ram[1205]=32'h1220000c; 
ram[1206]=32'h00000000; 
ram[1207]=32'h240400ff; 
ram[1208]=32'h1612fff7; 
ram[1209]=32'h00000000; 
ram[1210]=32'h0fc005fd; 
ram[1211]=32'h00000000; 
ram[1212]=32'h240400ff; 
ram[1213]=32'h00008021; 
ram[1214]=32'h0fc005e9; 
ram[1215]=32'h00000000; 
ram[1216]=32'h0bc0047d; 
ram[1217]=32'h00000000; 
ram[1218]=32'h0fc005fd; 
ram[1219]=32'h00000000; 
ram[1220]=32'h240400ff; 
ram[1221]=32'h0fc005e9; 
ram[1222]=32'h00000000; 
ram[1223]=32'h0bc0047d; 
ram[1224]=32'h00000000; 
ram[1225]=32'h27bdffd0; 
ram[1226]=32'hafb1001c; 
ram[1227]=32'h00808821; 
ram[1228]=32'h00002021; 
ram[1229]=32'hafbf002c; 
ram[1230]=32'hafb40028; 
ram[1231]=32'hafb20020; 
ram[1232]=32'hafb00018; 
ram[1233]=32'h30b400ff; 
ram[1234]=32'h00c08021; 
ram[1235]=32'hafb30024; 
ram[1236]=32'h0fc005f5; 
ram[1237]=32'h00000000; 
ram[1238]=32'h24040019; 
ram[1239]=32'h00112a40; 
ram[1240]=32'h240600ff; 
ram[1241]=32'h0fc002be; 
ram[1242]=32'h00000000; 
ram[1243]=32'h00409021; 
ram[1244]=32'h14400062; 
ram[1245]=32'h00000000; 
ram[1246]=32'h00009821; 
ram[1247]=32'h24110005; 
ram[1248]=32'h2631ffff; 
ram[1249]=32'h240400ff; 
ram[1250]=32'h3231ffff; 
ram[1251]=32'h0fc005e9; 
ram[1252]=32'h00000000; 
ram[1253]=32'h1620fffa; 
ram[1254]=32'h00000000; 
ram[1255]=32'h240400fc; 
ram[1256]=32'h26110200; 
ram[1257]=32'h0fc005e9; 
ram[1258]=32'h00000000; 
ram[1259]=32'h26100001; 
ram[1260]=32'h9204ffff; 
ram[1261]=32'h0fc005e9; 
ram[1262]=32'h00000000; 
ram[1263]=32'h1611fffb; 
ram[1264]=32'h00000000; 
ram[1265]=32'h240400ff; 
ram[1266]=32'h0fc005e9; 
ram[1267]=32'h00000000; 
ram[1268]=32'h26730001; 
ram[1269]=32'h240400ff; 
ram[1270]=32'h3273ffff; 
ram[1271]=32'h0fc005e9; 
ram[1272]=32'h00000000; 
ram[1273]=32'h240400ff; 
ram[1274]=32'h0fc005e9; 
ram[1275]=32'h00000000; 
ram[1276]=32'h2e6300ff; 
ram[1277]=32'h00409021; 
ram[1278]=32'h10600040; 
ram[1279]=32'h00000000; 
ram[1280]=32'h3052001f; 
ram[1281]=32'h24020005; 
ram[1282]=32'h1642ffdc; 
ram[1283]=32'h00000000; 
ram[1284]=32'h240400ff; 
ram[1285]=32'h0fc005e9; 
ram[1286]=32'h00000000; 
ram[1287]=32'h00409021; 
ram[1288]=32'h24117530; 
ram[1289]=32'h241300ff; 
ram[1290]=32'h0bc00513; 
ram[1291]=32'h00000000; 
ram[1292]=32'h2631ffff; 
ram[1293]=32'h0fc005e9; 
ram[1294]=32'h00000000; 
ram[1295]=32'h3231ffff; 
ram[1296]=32'h00409021; 
ram[1297]=32'h1220002d; 
ram[1298]=32'h00000000; 
ram[1299]=32'h240400ff; 
ram[1300]=32'h1653fff7; 
ram[1301]=32'h00000000; 
ram[1302]=32'h2694ffff; 
ram[1303]=32'h329400ff; 
ram[1304]=32'h1680ffc5; 
ram[1305]=32'h00000000; 
ram[1306]=32'h240400fd; 
ram[1307]=32'h0fc005e9; 
ram[1308]=32'h00000000; 
ram[1309]=32'h240400ff; 
ram[1310]=32'h0fc005e9; 
ram[1311]=32'h00000000; 
ram[1312]=32'h00409021; 
ram[1313]=32'h24107530; 
ram[1314]=32'h241100ff; 
ram[1315]=32'h0bc0052c; 
ram[1316]=32'h00000000; 
ram[1317]=32'h2610ffff; 
ram[1318]=32'h0fc005e9; 
ram[1319]=32'h00000000; 
ram[1320]=32'h3210ffff; 
ram[1321]=32'h00409021; 
ram[1322]=32'h12000014; 
ram[1323]=32'h00000000; 
ram[1324]=32'h240400ff; 
ram[1325]=32'h1651fff7; 
ram[1326]=32'h00000000; 
ram[1327]=32'h0fc005fd; 
ram[1328]=32'h00000000; 
ram[1329]=32'h240400ff; 
ram[1330]=32'h0fc005e9; 
ram[1331]=32'h00000000; 
ram[1332]=32'h8fbf002c; 
ram[1333]=32'h00009021; 
ram[1334]=32'h02401021; 
ram[1335]=32'h8fb40028; 
ram[1336]=32'h8fb30024; 
ram[1337]=32'h8fb20020; 
ram[1338]=32'h8fb1001c; 
ram[1339]=32'h8fb00018; 
ram[1340]=32'h27bd0030; 
ram[1341]=32'h03e00008; 
ram[1342]=32'h00000000; 
ram[1343]=32'h0fc005fd; 
ram[1344]=32'h00000000; 
ram[1345]=32'h240400ff; 
ram[1346]=32'h0fc005e9; 
ram[1347]=32'h00000000; 
ram[1348]=32'h8fbf002c; 
ram[1349]=32'h02401021; 
ram[1350]=32'h8fb40028; 
ram[1351]=32'h8fb30024; 
ram[1352]=32'h8fb20020; 
ram[1353]=32'h8fb1001c; 
ram[1354]=32'h8fb00018; 
ram[1355]=32'h27bd0030; 
ram[1356]=32'h03e00008; 
ram[1357]=32'h00000000; 
ram[1358]=32'h27bdffd8; 
ram[1359]=32'hafb1001c; 
ram[1360]=32'h00808821; 
ram[1361]=32'h00002021; 
ram[1362]=32'hafbf0024; 
ram[1363]=32'hafb00018; 
ram[1364]=32'hafb20020; 
ram[1365]=32'h0fc005f5; 
ram[1366]=32'h00000000; 
ram[1367]=32'h24040009; 
ram[1368]=32'h00002821; 
ram[1369]=32'h240600ff; 
ram[1370]=32'h241000fe; 
ram[1371]=32'h0fc002be; 
ram[1372]=32'h00000000; 
ram[1373]=32'h0bc00565; 
ram[1374]=32'h00000000; 
ram[1375]=32'h2610ffff; 
ram[1376]=32'h3210ffff; 
ram[1377]=32'h0fc002be; 
ram[1378]=32'h00000000; 
ram[1379]=32'h12000031; 
ram[1380]=32'h00000000; 
ram[1381]=32'h24040009; 
ram[1382]=32'h00002821; 
ram[1383]=32'h240600ff; 
ram[1384]=32'h1440fff6; 
ram[1385]=32'h00000000; 
ram[1386]=32'h240400ff; 
ram[1387]=32'h0fc005e9; 
ram[1388]=32'h00000000; 
ram[1389]=32'h24107530; 
ram[1390]=32'h241200fe; 
ram[1391]=32'h0bc00577; 
ram[1392]=32'h00000000; 
ram[1393]=32'h2610ffff; 
ram[1394]=32'h3210ffff; 
ram[1395]=32'h0fc005e9; 
ram[1396]=32'h00000000; 
ram[1397]=32'h1200001f; 
ram[1398]=32'h00000000; 
ram[1399]=32'h240400ff; 
ram[1400]=32'h1452fff8; 
ram[1401]=32'h00000000; 
ram[1402]=32'h26300010; 
ram[1403]=32'h240400ff; 
ram[1404]=32'h0fc005e9; 
ram[1405]=32'h00000000; 
ram[1406]=32'h26310001; 
ram[1407]=32'ha222ffff; 
ram[1408]=32'h1630fffa; 
ram[1409]=32'h00000000; 
ram[1410]=32'h240400ff; 
ram[1411]=32'h0fc005e9; 
ram[1412]=32'h00000000; 
ram[1413]=32'h240400ff; 
ram[1414]=32'h0fc005e9; 
ram[1415]=32'h00000000; 
ram[1416]=32'h0fc005fd; 
ram[1417]=32'h00000000; 
ram[1418]=32'h240400ff; 
ram[1419]=32'h0fc005e9; 
ram[1420]=32'h00000000; 
ram[1421]=32'h8fbf0024; 
ram[1422]=32'h8fb20020; 
ram[1423]=32'h8fb1001c; 
ram[1424]=32'h8fb00018; 
ram[1425]=32'h00001021; 
ram[1426]=32'h27bd0028; 
ram[1427]=32'h03e00008; 
ram[1428]=32'h00000000; 
ram[1429]=32'h0fc005fd; 
ram[1430]=32'h00000000; 
ram[1431]=32'h240400ff; 
ram[1432]=32'h0fc005e9; 
ram[1433]=32'h00000000; 
ram[1434]=32'h8fbf0024; 
ram[1435]=32'h8fb20020; 
ram[1436]=32'h8fb1001c; 
ram[1437]=32'h8fb00018; 
ram[1438]=32'h240200ff; 
ram[1439]=32'h27bd0028; 
ram[1440]=32'h03e00008; 
ram[1441]=32'h00000000; 
ram[1442]=32'h27bdffd0; 
ram[1443]=32'h27a40018; 
ram[1444]=32'hafbf002c; 
ram[1445]=32'h0fc0054e; 
ram[1446]=32'h00000000; 
ram[1447]=32'h8fa20018; 
ram[1448]=32'h304200c0; 
ram[1449]=32'h10400017; 
ram[1450]=32'h00000000; 
ram[1451]=32'h24030040; 
ram[1452]=32'h10430006; 
ram[1453]=32'h00000000; 
ram[1454]=32'h8fbf002c; 
ram[1455]=32'h00001021; 
ram[1456]=32'h27bd0030; 
ram[1457]=32'h03e00008; 
ram[1458]=32'h00000000; 
ram[1459]=32'h8fa2001c; 
ram[1460]=32'h93a40021; 
ram[1461]=32'h93a30020; 
ram[1462]=32'h00021682; 
ram[1463]=32'h00021400; 
ram[1464]=32'h00441025; 
ram[1465]=32'h00031a00; 
ram[1466]=32'h8fbf002c; 
ram[1467]=32'h00431025; 
ram[1468]=32'h24420001; 
ram[1469]=32'h00021280; 
ram[1470]=32'h27bd0030; 
ram[1471]=32'h03e00008; 
ram[1472]=32'h00000000; 
ram[1473]=32'h8fa30020; 
ram[1474]=32'h8fa4001c; 
ram[1475]=32'h93a2001f; 
ram[1476]=32'h00043182; 
ram[1477]=32'h000339c2; 
ram[1478]=32'h00032dc2; 
ram[1479]=32'h00021080; 
ram[1480]=32'h00031982; 
ram[1481]=32'h30e70006; 
ram[1482]=32'h30c60c00; 
ram[1483]=32'h30a50001; 
ram[1484]=32'h00042202; 
ram[1485]=32'h00c23025; 
ram[1486]=32'h00e52825; 
ram[1487]=32'h30620003; 
ram[1488]=32'h3084000f; 
ram[1489]=32'h8fbf002c; 
ram[1490]=32'h00461025; 
ram[1491]=32'h00a42021; 
ram[1492]=32'h24840002; 
ram[1493]=32'h24420001; 
ram[1494]=32'h00821004; 
ram[1495]=32'h27bd0030; 
ram[1496]=32'h03e00008; 
ram[1497]=32'h00000000; 
ram[1498]=32'h00000000; 
ram[1499]=32'h00000000; 
ram[1500]=32'h3c02b800; 
ram[1501]=32'h24030050; 
ram[1502]=32'ha0430500; 
ram[1503]=32'h24030002; 
ram[1504]=32'ha043050c; 
ram[1505]=32'h03e00008; 
ram[1506]=32'h00000000; 
ram[1507]=32'h3c02b800; 
ram[1508]=32'h90420504; 
ram[1509]=32'h30420001; 
ram[1510]=32'h38420001; 
ram[1511]=32'h03e00008; 
ram[1512]=32'h00000000; 
ram[1513]=32'h308400ff; 
ram[1514]=32'h3c02b800; 
ram[1515]=32'ha0440508; 
ram[1516]=32'h3c02b800; 
ram[1517]=32'h90430504; 
ram[1518]=32'h30630001; 
ram[1519]=32'h1460fffc; 
ram[1520]=32'h00000000; 
ram[1521]=32'h90420508; 
ram[1522]=32'h304200ff; 
ram[1523]=32'h03e00008; 
ram[1524]=32'h00000000; 
ram[1525]=32'h24020001; 
ram[1526]=32'h00822004; 
ram[1527]=32'h00041027; 
ram[1528]=32'h304200ff; 
ram[1529]=32'h3c03b800; 
ram[1530]=32'ha0620510; 
ram[1531]=32'h03e00008; 
ram[1532]=32'h00000000; 
ram[1533]=32'h2403000f; 
ram[1534]=32'h3c02b800; 
ram[1535]=32'ha0430510; 
ram[1536]=32'h03e00008; 
ram[1537]=32'h00000000; 
ram[1538]=32'h00000000; 
ram[1539]=32'h00000000; 
ram[1540]=32'h80820000; 
ram[1541]=32'h10400009; 
ram[1542]=32'h00000000; 
ram[1543]=32'h00801021; 
ram[1544]=32'h24420001; 
ram[1545]=32'h80430000; 
ram[1546]=32'h1460fffd; 
ram[1547]=32'h00000000; 
ram[1548]=32'h00441023; 
ram[1549]=32'h03e00008; 
ram[1550]=32'h00000000; 
ram[1551]=32'h00001021; 
ram[1552]=32'h03e00008; 
ram[1553]=32'h00000000; 
ram[1554]=32'h80a30000; 
ram[1555]=32'h00801021; 
ram[1556]=32'h00803021; 
ram[1557]=32'h10600007; 
ram[1558]=32'h00000000; 
ram[1559]=32'h24c60001; 
ram[1560]=32'h24a50001; 
ram[1561]=32'ha0c3ffff; 
ram[1562]=32'h80a30000; 
ram[1563]=32'h1460fffb; 
ram[1564]=32'h00000000; 
ram[1565]=32'ha0c00000; 
ram[1566]=32'h03e00008; 
ram[1567]=32'h00000000; 
ram[1568]=32'h80830000; 
ram[1569]=32'h00801021; 
ram[1570]=32'h10600014; 
ram[1571]=32'h00000000; 
ram[1572]=32'h00801821; 
ram[1573]=32'h24630001; 
ram[1574]=32'h80660000; 
ram[1575]=32'h14c0fffd; 
ram[1576]=32'h00000000; 
ram[1577]=32'h00621823; 
ram[1578]=32'h80a60000; 
ram[1579]=32'h00431821; 
ram[1580]=32'h10c00007; 
ram[1581]=32'h00000000; 
ram[1582]=32'h24630001; 
ram[1583]=32'h24a50001; 
ram[1584]=32'ha066ffff; 
ram[1585]=32'h80a60000; 
ram[1586]=32'h14c0fffb; 
ram[1587]=32'h00000000; 
ram[1588]=32'ha0600000; 
ram[1589]=32'h03e00008; 
ram[1590]=32'h00000000; 
ram[1591]=32'h00001821; 
ram[1592]=32'h0bc0062a; 
ram[1593]=32'h00000000; 
ram[1594]=32'h80a30000; 
ram[1595]=32'h00801021; 
ram[1596]=32'h10600012; 
ram[1597]=32'h00000000; 
ram[1598]=32'h18c00010; 
ram[1599]=32'h00000000; 
ram[1600]=32'h00a63021; 
ram[1601]=32'h00803821; 
ram[1602]=32'h0bc00646; 
ram[1603]=32'h00000000; 
ram[1604]=32'h10a60007; 
ram[1605]=32'h00000000; 
ram[1606]=32'h24e70001; 
ram[1607]=32'h24a50001; 
ram[1608]=32'ha0e3ffff; 
ram[1609]=32'h80a30000; 
ram[1610]=32'h1460fff9; 
ram[1611]=32'h00000000; 
ram[1612]=32'ha0e00000; 
ram[1613]=32'h03e00008; 
ram[1614]=32'h00000000; 
ram[1615]=32'h00403821; 
ram[1616]=32'h0bc0064c; 
ram[1617]=32'h00000000; 
ram[1618]=32'h80830000; 
ram[1619]=32'h00801021; 
ram[1620]=32'h1060001b; 
ram[1621]=32'h00000000; 
ram[1622]=32'h00801821; 
ram[1623]=32'h24630001; 
ram[1624]=32'h80670000; 
ram[1625]=32'h14e0fffd; 
ram[1626]=32'h00000000; 
ram[1627]=32'h00621823; 
ram[1628]=32'h80a70000; 
ram[1629]=32'h00431821; 
ram[1630]=32'h10e0000e; 
ram[1631]=32'h00000000; 
ram[1632]=32'h18c0000c; 
ram[1633]=32'h00000000; 
ram[1634]=32'h00a63021; 
ram[1635]=32'h0bc00667; 
ram[1636]=32'h00000000; 
ram[1637]=32'h10a60007; 
ram[1638]=32'h00000000; 
ram[1639]=32'h24630001; 
ram[1640]=32'h24a50001; 
ram[1641]=32'ha067ffff; 
ram[1642]=32'h80a70000; 
ram[1643]=32'h14e0fff9; 
ram[1644]=32'h00000000; 
ram[1645]=32'ha0600000; 
ram[1646]=32'h03e00008; 
ram[1647]=32'h00000000; 
ram[1648]=32'h00001821; 
ram[1649]=32'h0bc0065c; 
ram[1650]=32'h00000000; 
ram[1651]=32'h0bc0067b; 
ram[1652]=32'h00000000; 
ram[1653]=32'h24a50001; 
ram[1654]=32'h00c31023; 
ram[1655]=32'h10600008; 
ram[1656]=32'h00000000; 
ram[1657]=32'h14400007; 
ram[1658]=32'h00000000; 
ram[1659]=32'h80860000; 
ram[1660]=32'h80a30000; 
ram[1661]=32'h24840001; 
ram[1662]=32'h14c0fff6; 
ram[1663]=32'h00000000; 
ram[1664]=32'h00c31023; 
ram[1665]=32'h03e00008; 
ram[1666]=32'h00000000; 
ram[1667]=32'h80830000; 
ram[1668]=32'h1060001b; 
ram[1669]=32'h00000000; 
ram[1670]=32'h80a20000; 
ram[1671]=32'h10400018; 
ram[1672]=32'h00000000; 
ram[1673]=32'h18c00016; 
ram[1674]=32'h00000000; 
ram[1675]=32'h00621023; 
ram[1676]=32'h24840001; 
ram[1677]=32'h24a50001; 
ram[1678]=32'h1040000d; 
ram[1679]=32'h00000000; 
ram[1680]=32'h0bc006a9; 
ram[1681]=32'h00000000; 
ram[1682]=32'h80a70000; 
ram[1683]=32'h24840001; 
ram[1684]=32'h00671023; 
ram[1685]=32'h10e0000a; 
ram[1686]=32'h00000000; 
ram[1687]=32'h10c0000e; 
ram[1688]=32'h00000000; 
ram[1689]=32'h24a50001; 
ram[1690]=32'h1440000c; 
ram[1691]=32'h00000000; 
ram[1692]=32'h80830000; 
ram[1693]=32'h24c6ffff; 
ram[1694]=32'h1460fff3; 
ram[1695]=32'h00000000; 
ram[1696]=32'h10c00005; 
ram[1697]=32'h00000000; 
ram[1698]=32'h80a20000; 
ram[1699]=32'h00621023; 
ram[1700]=32'h03e00008; 
ram[1701]=32'h00000000; 
ram[1702]=32'h00001021; 
ram[1703]=32'h03e00008; 
ram[1704]=32'h00000000; 
ram[1705]=32'h03e00008; 
ram[1706]=32'h00000000; 
ram[1707]=32'h00801021; 
ram[1708]=32'h10c00009; 
ram[1709]=32'h00000000; 
ram[1710]=32'h00a63021; 
ram[1711]=32'h00801821; 
ram[1712]=32'h24a50001; 
ram[1713]=32'h90a7ffff; 
ram[1714]=32'h24630001; 
ram[1715]=32'ha067ffff; 
ram[1716]=32'h14a6fffb; 
ram[1717]=32'h00000000; 
ram[1718]=32'h03e00008; 
ram[1719]=32'h00000000; 
ram[1720]=32'h00801021; 
ram[1721]=32'h24c7ffff; 
ram[1722]=32'h00801821; 
ram[1723]=32'h2408ffff; 
ram[1724]=32'h10c00008; 
ram[1725]=32'h00000000; 
ram[1726]=32'h24a50004; 
ram[1727]=32'h8ca6fffc; 
ram[1728]=32'h24630004; 
ram[1729]=32'h24e7ffff; 
ram[1730]=32'hac66fffc; 
ram[1731]=32'h14e8fffa; 
ram[1732]=32'h00000000; 
ram[1733]=32'h03e00008; 
ram[1734]=32'h00000000; 
ram[1735]=32'h00801021; 
ram[1736]=32'h30a500ff; 
ram[1737]=32'h10c00007; 
ram[1738]=32'h00000000; 
ram[1739]=32'h00863021; 
ram[1740]=32'h00801821; 
ram[1741]=32'h24630001; 
ram[1742]=32'ha065ffff; 
ram[1743]=32'h1466fffd; 
ram[1744]=32'h00000000; 
ram[1745]=32'h03e00008; 
ram[1746]=32'h00000000; 
ram[1747]=32'h00801021; 
ram[1748]=32'h30a5ffff; 
ram[1749]=32'h24c7ffff; 
ram[1750]=32'h00801821; 
ram[1751]=32'h2408ffff; 
ram[1752]=32'h10c00006; 
ram[1753]=32'h00000000; 
ram[1754]=32'h24630002; 
ram[1755]=32'h24e7ffff; 
ram[1756]=32'ha465fffe; 
ram[1757]=32'h14e8fffc; 
ram[1758]=32'h00000000; 
ram[1759]=32'h03e00008; 
ram[1760]=32'h00000000; 
ram[1761]=32'h18c00011; 
ram[1762]=32'h00000000; 
ram[1763]=32'h80870000; 
ram[1764]=32'h80a20000; 
ram[1765]=32'h00001821; 
ram[1766]=32'h10e20007; 
ram[1767]=32'h00000000; 
ram[1768]=32'h0bc006f6; 
ram[1769]=32'h00000000; 
ram[1770]=32'h80e70000; 
ram[1771]=32'h80420000; 
ram[1772]=32'h14e20009; 
ram[1773]=32'h00000000; 
ram[1774]=32'h24630001; 
ram[1775]=32'h00833821; 
ram[1776]=32'h00a31021; 
ram[1777]=32'h1466fff8; 
ram[1778]=32'h00000000; 
ram[1779]=32'h00001021; 
ram[1780]=32'h03e00008; 
ram[1781]=32'h00000000; 
ram[1782]=32'h00e21023; 
ram[1783]=32'h03e00008; 
ram[1784]=32'h00000000; 
ram[1785]=32'haca00000; 
ram[1786]=32'h80820000; 
ram[1787]=32'h10400018; 
ram[1788]=32'h00000000; 
ram[1789]=32'h2443ffd0; 
ram[1790]=32'h306300ff; 
ram[1791]=32'h2c63000a; 
ram[1792]=32'h10600016; 
ram[1793]=32'h00000000; 
ram[1794]=32'h00001821; 
ram[1795]=32'h0bc00707; 
ram[1796]=32'h00000000; 
ram[1797]=32'h10c00011; 
ram[1798]=32'h00000000; 
ram[1799]=32'h00033040; 
ram[1800]=32'h000318c0; 
ram[1801]=32'h00c31821; 
ram[1802]=32'h00621021; 
ram[1803]=32'h2443ffd0; 
ram[1804]=32'haca30000; 
ram[1805]=32'h24840001; 
ram[1806]=32'h80820000; 
ram[1807]=32'h2446ffd0; 
ram[1808]=32'h30c600ff; 
ram[1809]=32'h2cc6000a; 
ram[1810]=32'h1440fff2; 
ram[1811]=32'h00000000; 
ram[1812]=32'h00001021; 
ram[1813]=32'h03e00008; 
ram[1814]=32'h00000000; 
ram[1815]=32'h2402ffff; 
ram[1816]=32'h03e00008; 
ram[1817]=32'h00000000; 
ram[1818]=32'h04800030; 
ram[1819]=32'h00000000; 
ram[1820]=32'h10800029; 
ram[1821]=32'h00000000; 
ram[1822]=32'h3c076666; 
ram[1823]=32'h00801021; 
ram[1824]=32'h00003021; 
ram[1825]=32'h24e76667; 
ram[1826]=32'h0bc00725; 
ram[1827]=32'h00000000; 
ram[1828]=32'h00603021; 
ram[1829]=32'h00470018; 
ram[1830]=32'h000217c3; 
ram[1831]=32'h00001810; 
ram[1832]=32'h00031883; 
ram[1833]=32'h00621023; 
ram[1834]=32'h24c30001; 
ram[1835]=32'h1440fff8; 
ram[1836]=32'h00000000; 
ram[1837]=32'h00a62821; 
ram[1838]=32'h3c096666; 
ram[1839]=32'ha0a00001; 
ram[1840]=32'h00a01021; 
ram[1841]=32'h25296667; 
ram[1842]=32'h00890018; 
ram[1843]=32'h00043fc3; 
ram[1844]=32'h00001810; 
ram[1845]=32'h2442ffff; 
ram[1846]=32'h00031883; 
ram[1847]=32'h00671823; 
ram[1848]=32'h000338c0; 
ram[1849]=32'h00034040; 
ram[1850]=32'h01074021; 
ram[1851]=32'h24470001; 
ram[1852]=32'h00882023; 
ram[1853]=32'h00e63821; 
ram[1854]=32'h24840030; 
ram[1855]=32'h00e53823; 
ram[1856]=32'ha0440001; 
ram[1857]=32'h00602021; 
ram[1858]=32'h1ce0ffef; 
ram[1859]=32'h00000000; 
ram[1860]=32'h03e00008; 
ram[1861]=32'h00000000; 
ram[1862]=32'h24020030; 
ram[1863]=32'ha0a20000; 
ram[1864]=32'ha0a00001; 
ram[1865]=32'h03e00008; 
ram[1866]=32'h00000000; 
ram[1867]=32'h2402002d; 
ram[1868]=32'ha0a20000; 
ram[1869]=32'h00042023; 
ram[1870]=32'h24a50001; 
ram[1871]=32'h0bc0071e; 
ram[1872]=32'h00000000; 
ram[1873]=32'h00000000; 
ram[1874]=32'h00000000; 
ram[1875]=32'h00000000; 
ram[1876]=32'h27bdff90; 
ram[1877]=32'hafb60060; 
ram[1878]=32'h3c169f00; 
ram[1879]=32'hafb70064; 
ram[1880]=32'hafb5005c; 
ram[1881]=32'hafb40058; 
ram[1882]=32'hafb00048; 
ram[1883]=32'hafbf006c; 
ram[1884]=32'hafbe0068; 
ram[1885]=32'hafb30054; 
ram[1886]=32'hafb20050; 
ram[1887]=32'hafb1004c; 
ram[1888]=32'hafa40038; 
ram[1889]=32'h00808021; 
ram[1890]=32'h24150025; 
ram[1891]=32'h24170063; 
ram[1892]=32'h27b40018; 
ram[1893]=32'h26d62930; 
ram[1894]=32'h80a30000; 
ram[1895]=32'h10600009; 
ram[1896]=32'h00000000; 
ram[1897]=32'h10750016; 
ram[1898]=32'h00000000; 
ram[1899]=32'ha2030000; 
ram[1900]=32'h24a50001; 
ram[1901]=32'h80a30000; 
ram[1902]=32'h26100001; 
ram[1903]=32'h1460fff9; 
ram[1904]=32'h00000000; 
ram[1905]=32'ha2000000; 
ram[1906]=32'h8fa40038; 
ram[1907]=32'h8fbf006c; 
ram[1908]=32'h8fbe0068; 
ram[1909]=32'h8fb70064; 
ram[1910]=32'h8fb60060; 
ram[1911]=32'h8fb5005c; 
ram[1912]=32'h8fb40058; 
ram[1913]=32'h8fb30054; 
ram[1914]=32'h8fb20050; 
ram[1915]=32'h8fb1004c; 
ram[1916]=32'h8fb00048; 
ram[1917]=32'h27bd0070; 
ram[1918]=32'h0bc00604; 
ram[1919]=32'h00000000; 
ram[1920]=32'h80a20001; 
ram[1921]=32'h24b10001; 
ram[1922]=32'h00009821; 
ram[1923]=32'h00009021; 
ram[1924]=32'h00005821; 
ram[1925]=32'h00005021; 
ram[1926]=32'h0000f021; 
ram[1927]=32'h240c0073; 
ram[1928]=32'h24190075; 
ram[1929]=32'h24180064; 
ram[1930]=32'h240e006f; 
ram[1931]=32'h2409002d; 
ram[1932]=32'h24040001; 
ram[1933]=32'h240d002e; 
ram[1934]=32'h240f0030; 
ram[1935]=32'h10570069; 
ram[1936]=32'h00000000; 
ram[1937]=32'h28470064; 
ram[1938]=32'h10e00010; 
ram[1939]=32'h00000000; 
ram[1940]=32'h10490086; 
ram[1941]=32'h00000000; 
ram[1942]=32'h2847002e; 
ram[1943]=32'h10e00058; 
ram[1944]=32'h00000000; 
ram[1945]=32'h10400073; 
ram[1946]=32'h00000000; 
ram[1947]=32'h145500af; 
ram[1948]=32'h00000000; 
ram[1949]=32'h26220001; 
ram[1950]=32'ha2150000; 
ram[1951]=32'h00402821; 
ram[1952]=32'h26100001; 
ram[1953]=32'h0bc00766; 
ram[1954]=32'h00000000; 
ram[1955]=32'h104c007e; 
ram[1956]=32'h00000000; 
ram[1957]=32'h28470074; 
ram[1958]=32'h10e0009f; 
ram[1959]=32'h00000000; 
ram[1960]=32'h10580003; 
ram[1961]=32'h00000000; 
ram[1962]=32'h144e00a0; 
ram[1963]=32'h00000000; 
ram[1964]=32'h8cc30000; 
ram[1965]=32'h24c60004; 
ram[1966]=32'h146000c7; 
ram[1967]=32'h00000000; 
ram[1968]=32'h24020030; 
ram[1969]=32'ha3a20018; 
ram[1970]=32'h24020001; 
ram[1971]=32'h0053202a; 
ram[1972]=32'h02603821; 
ram[1973]=32'h00006021; 
ram[1974]=32'h24030001; 
ram[1975]=32'ha3a00019; 
ram[1976]=32'h24050030; 
ram[1977]=32'h24090001; 
ram[1978]=32'h000b500b; 
ram[1979]=32'h0044380a; 
ram[1980]=32'h118300dc; 
ram[1981]=32'h00000000; 
ram[1982]=32'h13c301b6; 
ram[1983]=32'h00000000; 
ram[1984]=32'h00f2182a; 
ram[1985]=32'h1060019a; 
ram[1986]=32'h00000000; 
ram[1987]=32'h02471823; 
ram[1988]=32'h24040030; 
ram[1989]=32'h24080020; 
ram[1990]=32'h02031821; 
ram[1991]=32'h010a200a; 
ram[1992]=32'h26100001; 
ram[1993]=32'ha204ffff; 
ram[1994]=32'h1603fffd; 
ram[1995]=32'h00000000; 
ram[1996]=32'h0047202a; 
ram[1997]=32'h10800174; 
ram[1998]=32'h00000000; 
ram[1999]=32'h00e28023; 
ram[2000]=32'h00708021; 
ram[2001]=32'h24020030; 
ram[2002]=32'h24630001; 
ram[2003]=32'ha062ffff; 
ram[2004]=32'h1470fffd; 
ram[2005]=32'h00000000; 
ram[2006]=32'h10a0016e; 
ram[2007]=32'h00000000; 
ram[2008]=32'h27a40019; 
ram[2009]=32'h00801821; 
ram[2010]=32'h24840001; 
ram[2011]=32'h8085ffff; 
ram[2012]=32'h14a0fffc; 
ram[2013]=32'h00000000; 
ram[2014]=32'h02002821; 
ram[2015]=32'h0bc007e2; 
ram[2016]=32'h00000000; 
ram[2017]=32'h00802821; 
ram[2018]=32'h2463ffff; 
ram[2019]=32'h90680000; 
ram[2020]=32'h0283382b; 
ram[2021]=32'h24a40001; 
ram[2022]=32'ha0a80000; 
ram[2023]=32'h14e0fff9; 
ram[2024]=32'h00000000; 
ram[2025]=32'h02098021; 
ram[2026]=32'ha0a00001; 
ram[2027]=32'h26220001; 
ram[2028]=32'ha2000000; 
ram[2029]=32'h00402821; 
ram[2030]=32'h0bc00766; 
ram[2031]=32'h00000000; 
ram[2032]=32'h104d006c; 
ram[2033]=32'h00000000; 
ram[2034]=32'h144f0058; 
ram[2035]=32'h00000000; 
ram[2036]=32'h82220001; 
ram[2037]=32'h240a0001; 
ram[2038]=32'h26310001; 
ram[2039]=32'h1457ff99; 
ram[2040]=32'h00000000; 
ram[2041]=32'h17c000b4; 
ram[2042]=32'h00000000; 
ram[2043]=32'h2a420002; 
ram[2044]=32'h14400142; 
ram[2045]=32'h00000000; 
ram[2046]=32'h2652ffff; 
ram[2047]=32'h02129021; 
ram[2048]=32'h24020020; 
ram[2049]=32'h26100001; 
ram[2050]=32'ha202ffff; 
ram[2051]=32'h1612fffd; 
ram[2052]=32'h00000000; 
ram[2053]=32'h80c20000; 
ram[2054]=32'h26500001; 
ram[2055]=32'ha2420000; 
ram[2056]=32'h26220001; 
ram[2057]=32'h24c60004; 
ram[2058]=32'h00402821; 
ram[2059]=32'h0bc00766; 
ram[2060]=32'h00000000; 
ram[2061]=32'h8fbf006c; 
ram[2062]=32'h8fbe0068; 
ram[2063]=32'h8fb70064; 
ram[2064]=32'h8fb60060; 
ram[2065]=32'h8fb5005c; 
ram[2066]=32'h8fb40058; 
ram[2067]=32'h8fb30054; 
ram[2068]=32'h8fb20050; 
ram[2069]=32'h8fb1004c; 
ram[2070]=32'h8fb00048; 
ram[2071]=32'h00001021; 
ram[2072]=32'h27bd0070; 
ram[2073]=32'h03e00008; 
ram[2074]=32'h00000000; 
ram[2075]=32'h13c4012c; 
ram[2076]=32'h00000000; 
ram[2077]=32'h82220001; 
ram[2078]=32'h241e0001; 
ram[2079]=32'h26310001; 
ram[2080]=32'h0bc0078f; 
ram[2081]=32'h00000000; 
ram[2082]=32'h8cc50000; 
ram[2083]=32'h24c60004; 
ram[2084]=32'h00a02021; 
ram[2085]=32'hafa6003c; 
ram[2086]=32'hafa50040; 
ram[2087]=32'h0fc00604; 
ram[2088]=32'h00000000; 
ram[2089]=32'h00403021; 
ram[2090]=32'h8fa50040; 
ram[2091]=32'h12600003; 
ram[2092]=32'h00000000; 
ram[2093]=32'h0262102a; 
ram[2094]=32'h0262300b; 
ram[2095]=32'h17c000ad; 
ram[2096]=32'h00000000; 
ram[2097]=32'h00d2102a; 
ram[2098]=32'h104000da; 
ram[2099]=32'h00000000; 
ram[2100]=32'h02469023; 
ram[2101]=32'h02129021; 
ram[2102]=32'h24030020; 
ram[2103]=32'h26100001; 
ram[2104]=32'ha203ffff; 
ram[2105]=32'h1612fffd; 
ram[2106]=32'h00000000; 
ram[2107]=32'h02402021; 
ram[2108]=32'hafa60040; 
ram[2109]=32'h0fc00612; 
ram[2110]=32'h00000000; 
ram[2111]=32'h8fa60040; 
ram[2112]=32'h26220001; 
ram[2113]=32'h02468021; 
ram[2114]=32'h8fa6003c; 
ram[2115]=32'h00402821; 
ram[2116]=32'h0bc00766; 
ram[2117]=32'h00000000; 
ram[2118]=32'h1059ff65; 
ram[2119]=32'h00000000; 
ram[2120]=32'h24070078; 
ram[2121]=32'h1047ff62; 
ram[2122]=32'h00000000; 
ram[2123]=32'h2447ffd0; 
ram[2124]=32'h30e200ff; 
ram[2125]=32'h2c42000a; 
ram[2126]=32'h104000f9; 
ram[2127]=32'h00000000; 
ram[2128]=32'h26310001; 
ram[2129]=32'h00124040; 
ram[2130]=32'h82220000; 
ram[2131]=32'h001290c0; 
ram[2132]=32'h01129021; 
ram[2133]=32'h00f29021; 
ram[2134]=32'h2447ffd0; 
ram[2135]=32'h30e800ff; 
ram[2136]=32'h2d08000a; 
ram[2137]=32'h1500fff6; 
ram[2138]=32'h00000000; 
ram[2139]=32'h0bc0078f; 
ram[2140]=32'h00000000; 
ram[2141]=32'h116400ea; 
ram[2142]=32'h00000000; 
ram[2143]=32'h82220001; 
ram[2144]=32'h10490061; 
ram[2145]=32'h00000000; 
ram[2146]=32'h2447ffd0; 
ram[2147]=32'h30e800ff; 
ram[2148]=32'h2d08000a; 
ram[2149]=32'h26310001; 
ram[2150]=32'h1100000c; 
ram[2151]=32'h00000000; 
ram[2152]=32'h26310001; 
ram[2153]=32'h00134040; 
ram[2154]=32'h82220000; 
ram[2155]=32'h001398c0; 
ram[2156]=32'h01139821; 
ram[2157]=32'h00f39821; 
ram[2158]=32'h2447ffd0; 
ram[2159]=32'h30e800ff; 
ram[2160]=32'h2d08000a; 
ram[2161]=32'h1500fff6; 
ram[2162]=32'h00000000; 
ram[2163]=32'h240b0001; 
ram[2164]=32'h0bc0078f; 
ram[2165]=32'h00000000; 
ram[2166]=32'h24040064; 
ram[2167]=32'h1044005b; 
ram[2168]=32'h00000000; 
ram[2169]=32'h24040075; 
ram[2170]=32'h1044005a; 
ram[2171]=32'h00000000; 
ram[2172]=32'h24040078; 
ram[2173]=32'h10440074; 
ram[2174]=32'h00000000; 
ram[2175]=32'h3842006f; 
ram[2176]=32'h24040008; 
ram[2177]=32'h0002200b; 
ram[2178]=32'h00006021; 
ram[2179]=32'h00001021; 
ram[2180]=32'h0064001b; 
ram[2181]=32'h24420001; 
ram[2182]=32'h02822821; 
ram[2183]=32'h00003810; 
ram[2184]=32'h00001812; 
ram[2185]=32'h02c73821; 
ram[2186]=32'h90e70000; 
ram[2187]=32'ha0a7ffff; 
ram[2188]=32'h1460fff7; 
ram[2189]=32'h00000000; 
ram[2190]=32'h00404821; 
ram[2191]=32'h02821821; 
ram[2192]=32'ha0600000; 
ram[2193]=32'h0053202a; 
ram[2194]=32'h02603821; 
ram[2195]=32'h24030001; 
ram[2196]=32'h83a50018; 
ram[2197]=32'h000b500b; 
ram[2198]=32'h0044380a; 
ram[2199]=32'h1583ff26; 
ram[2200]=32'h00000000; 
ram[2201]=32'h24e80001; 
ram[2202]=32'h13cc0075; 
ram[2203]=32'h00000000; 
ram[2204]=32'h114c0059; 
ram[2205]=32'h00000000; 
ram[2206]=32'h0112182a; 
ram[2207]=32'h02002021; 
ram[2208]=32'h10600008; 
ram[2209]=32'h00000000; 
ram[2210]=32'h02482023; 
ram[2211]=32'h02042021; 
ram[2212]=32'h24030020; 
ram[2213]=32'h26100001; 
ram[2214]=32'ha203ffff; 
ram[2215]=32'h1604fffd; 
ram[2216]=32'h00000000; 
ram[2217]=32'h2408002d; 
ram[2218]=32'h24830001; 
ram[2219]=32'ha0880000; 
ram[2220]=32'h0bc007cc; 
ram[2221]=32'h00000000; 
ram[2222]=32'h80c30000; 
ram[2223]=32'h2a420002; 
ram[2224]=32'h26040001; 
ram[2225]=32'h24c60004; 
ram[2226]=32'ha2030000; 
ram[2227]=32'h144000b6; 
ram[2228]=32'h00000000; 
ram[2229]=32'h02128021; 
ram[2230]=32'h00801021; 
ram[2231]=32'h24030020; 
ram[2232]=32'h24420001; 
ram[2233]=32'ha043ffff; 
ram[2234]=32'h1450fffd; 
ram[2235]=32'h00000000; 
ram[2236]=32'h2650ffff; 
ram[2237]=32'h26220001; 
ram[2238]=32'h00908021; 
ram[2239]=32'h00402821; 
ram[2240]=32'h0bc00766; 
ram[2241]=32'h00000000; 
ram[2242]=32'h82220002; 
ram[2243]=32'h26310002; 
ram[2244]=32'h2447ffd0; 
ram[2245]=32'h30e700ff; 
ram[2246]=32'h2ce7000a; 
ram[2247]=32'h10e0ffab; 
ram[2248]=32'h00000000; 
ram[2249]=32'h26310001; 
ram[2250]=32'h82220000; 
ram[2251]=32'h2447ffd0; 
ram[2252]=32'h30e700ff; 
ram[2253]=32'h2ce7000a; 
ram[2254]=32'h14e0fffa; 
ram[2255]=32'h00000000; 
ram[2256]=32'h240b0001; 
ram[2257]=32'h0bc0078f; 
ram[2258]=32'h00000000; 
ram[2259]=32'h04600035; 
ram[2260]=32'h00000000; 
ram[2261]=32'h00006021; 
ram[2262]=32'h2404000a; 
ram[2263]=32'h1460ffab; 
ram[2264]=32'h00000000; 
ram[2265]=32'h00004821; 
ram[2266]=32'h00001021; 
ram[2267]=32'h0bc0088f; 
ram[2268]=32'h00000000; 
ram[2269]=32'h02002021; 
ram[2270]=32'hafa60040; 
ram[2271]=32'h0fc00612; 
ram[2272]=32'h00000000; 
ram[2273]=32'h8fa60040; 
ram[2274]=32'h00d2182a; 
ram[2275]=32'h02061021; 
ram[2276]=32'h1060008a; 
ram[2277]=32'h00000000; 
ram[2278]=32'h02463023; 
ram[2279]=32'h00468021; 
ram[2280]=32'h24030020; 
ram[2281]=32'h24420001; 
ram[2282]=32'ha043ffff; 
ram[2283]=32'h1450fffd; 
ram[2284]=32'h00000000; 
ram[2285]=32'h8fa6003c; 
ram[2286]=32'h26220001; 
ram[2287]=32'h00402821; 
ram[2288]=32'h0bc00766; 
ram[2289]=32'h00000000; 
ram[2290]=32'h24040010; 
ram[2291]=32'h00006021; 
ram[2292]=32'h0bc00883; 
ram[2293]=32'h00000000; 
ram[2294]=32'h240a002d; 
ram[2295]=32'h0112202a; 
ram[2296]=32'h26030001; 
ram[2297]=32'ha20a0000; 
ram[2298]=32'h1080fed1; 
ram[2299]=32'h00000000; 
ram[2300]=32'h26440001; 
ram[2301]=32'h00882023; 
ram[2302]=32'h02048021; 
ram[2303]=32'h240a0030; 
ram[2304]=32'h00602021; 
ram[2305]=32'h24840001; 
ram[2306]=32'ha08affff; 
ram[2307]=32'h1490fffd; 
ram[2308]=32'h00000000; 
ram[2309]=32'h02484023; 
ram[2310]=32'h00681821; 
ram[2311]=32'h0bc007cc; 
ram[2312]=32'h00000000; 
ram[2313]=32'h00031823; 
ram[2314]=32'h240c0001; 
ram[2315]=32'h0bc008d6; 
ram[2316]=32'h00000000; 
ram[2317]=32'h02009021; 
ram[2318]=32'h0bc0083b; 
ram[2319]=32'h00000000; 
ram[2320]=32'h2407002d; 
ram[2321]=32'h26030001; 
ram[2322]=32'ha2070000; 
ram[2323]=32'h10800053; 
ram[2324]=32'h00000000; 
ram[2325]=32'h02621023; 
ram[2326]=32'h00625021; 
ram[2327]=32'h24020030; 
ram[2328]=32'h24630001; 
ram[2329]=32'ha062ffff; 
ram[2330]=32'h146afffd; 
ram[2331]=32'h00000000; 
ram[2332]=32'h10a00047; 
ram[2333]=32'h00000000; 
ram[2334]=32'h27a30019; 
ram[2335]=32'h00601021; 
ram[2336]=32'h24630001; 
ram[2337]=32'h8064ffff; 
ram[2338]=32'h1480fffc; 
ram[2339]=32'h00000000; 
ram[2340]=32'h01402021; 
ram[2341]=32'h0bc00928; 
ram[2342]=32'h00000000; 
ram[2343]=32'h00602021; 
ram[2344]=32'h2442ffff; 
ram[2345]=32'h90470000; 
ram[2346]=32'h0282282b; 
ram[2347]=32'h24830001; 
ram[2348]=32'ha0870000; 
ram[2349]=32'h14a0fff9; 
ram[2350]=32'h00000000; 
ram[2351]=32'h0112182a; 
ram[2352]=32'ha0800001; 
ram[2353]=32'h01491021; 
ram[2354]=32'h1060002c; 
ram[2355]=32'h00000000; 
ram[2356]=32'h02484023; 
ram[2357]=32'h00488021; 
ram[2358]=32'h24030020; 
ram[2359]=32'h24420001; 
ram[2360]=32'ha043ffff; 
ram[2361]=32'h1450fffd; 
ram[2362]=32'h00000000; 
ram[2363]=32'ha2000000; 
ram[2364]=32'h26220001; 
ram[2365]=32'h0bc007ed; 
ram[2366]=32'h00000000; 
ram[2367]=32'h02009021; 
ram[2368]=32'h0bc00805; 
ram[2369]=32'h00000000; 
ram[2370]=32'h00608021; 
ram[2371]=32'h0bc007d6; 
ram[2372]=32'h00000000; 
ram[2373]=32'h02801821; 
ram[2374]=32'h0bc007de; 
ram[2375]=32'h00000000; 
ram[2376]=32'h0225102b; 
ram[2377]=32'h1440ffa4; 
ram[2378]=32'h00000000; 
ram[2379]=32'h26220001; 
ram[2380]=32'h02003821; 
ram[2381]=32'h00a02021; 
ram[2382]=32'h0bc00951; 
ram[2383]=32'h00000000; 
ram[2384]=32'h80830000; 
ram[2385]=32'h24e70001; 
ram[2386]=32'h24840001; 
ram[2387]=32'ha0e3ffff; 
ram[2388]=32'h1482fffb; 
ram[2389]=32'h00000000; 
ram[2390]=32'h02251823; 
ram[2391]=32'h24630001; 
ram[2392]=32'h02038021; 
ram[2393]=32'h00402821; 
ram[2394]=32'h0bc00766; 
ram[2395]=32'h00000000; 
ram[2396]=32'h02001821; 
ram[2397]=32'h0bc007cc; 
ram[2398]=32'h00000000; 
ram[2399]=32'h00408021; 
ram[2400]=32'ha2000000; 
ram[2401]=32'h26220001; 
ram[2402]=32'h0bc007ed; 
ram[2403]=32'h00000000; 
ram[2404]=32'h02801021; 
ram[2405]=32'h0bc00924; 
ram[2406]=32'h00000000; 
ram[2407]=32'h00605021; 
ram[2408]=32'h0bc0091c; 
ram[2409]=32'h00000000; 
ram[2410]=32'h26220001; 
ram[2411]=32'h00808021; 
ram[2412]=32'h00402821; 
ram[2413]=32'h0bc00766; 
ram[2414]=32'h00000000; 
ram[2415]=32'h00408021; 
ram[2416]=32'h26220001; 
ram[2417]=32'h8fa6003c; 
ram[2418]=32'h00402821; 
ram[2419]=32'h0bc00766; 
ram[2420]=32'h00000000; 
ram[2421]=32'h00e04021; 
ram[2422]=32'h02001821; 
ram[2423]=32'h0bc00913; 
ram[2424]=32'h00000000; 
ram[2425]=32'h27bdfbd8; 
ram[2426]=32'h00801821; 
ram[2427]=32'h00a01021; 
ram[2428]=32'h27a40018; 
ram[2429]=32'hafb1041c; 
ram[2430]=32'h00602821; 
ram[2431]=32'h00c08821; 
ram[2432]=32'h00403021; 
ram[2433]=32'hafb20420; 
ram[2434]=32'hafb00418; 
ram[2435]=32'hafbf0424; 
ram[2436]=32'h0fc00754; 
ram[2437]=32'h00000000; 
ram[2438]=32'h83a40018; 
ram[2439]=32'h00409021; 
ram[2440]=32'h27b00019; 
ram[2441]=32'h10800008; 
ram[2442]=32'h00000000; 
ram[2443]=32'h26100001; 
ram[2444]=32'h0220c821; 
ram[2445]=32'h0320f809; 
ram[2446]=32'h00000000; 
ram[2447]=32'h8204ffff; 
ram[2448]=32'h1480fffa; 
ram[2449]=32'h00000000; 
ram[2450]=32'h8fbf0424; 
ram[2451]=32'h02401021; 
ram[2452]=32'h8fb1041c; 
ram[2453]=32'h8fb20420; 
ram[2454]=32'h8fb00418; 
ram[2455]=32'h27bd0428; 
ram[2456]=32'h03e00008; 
ram[2457]=32'h00000000; 
ram[2458]=32'h27bdffe0; 
ram[2459]=32'hafa60028; 
ram[2460]=32'h27a60028; 
ram[2461]=32'hafbf001c; 
ram[2462]=32'hafa7002c; 
ram[2463]=32'hafa50024; 
ram[2464]=32'h0fc00754; 
ram[2465]=32'h00000000; 
ram[2466]=32'h8fbf001c; 
ram[2467]=32'h27bd0020; 
ram[2468]=32'h03e00008; 
ram[2469]=32'h00000000; 
ram[2470]=32'h80a20000; 
ram[2471]=32'h10400018; 
ram[2472]=32'h00000000; 
ram[2473]=32'h00a01021; 
ram[2474]=32'h24420001; 
ram[2475]=32'h80430000; 
ram[2476]=32'h1460fffd; 
ram[2477]=32'h00000000; 
ram[2478]=32'h2442ffff; 
ram[2479]=32'h80470000; 
ram[2480]=32'h00a2302b; 
ram[2481]=32'h24830001; 
ram[2482]=32'ha0870000; 
ram[2483]=32'h10c00009; 
ram[2484]=32'h00000000; 
ram[2485]=32'h00602021; 
ram[2486]=32'h2442ffff; 
ram[2487]=32'h80470000; 
ram[2488]=32'h00a2302b; 
ram[2489]=32'h24830001; 
ram[2490]=32'ha0870000; 
ram[2491]=32'h14c0fff9; 
ram[2492]=32'h00000000; 
ram[2493]=32'ha0800001; 
ram[2494]=32'h03e00008; 
ram[2495]=32'h00000000; 
ram[2496]=32'h00a01021; 
ram[2497]=32'h0bc009b6; 
ram[2498]=32'h00000000; 
ram[2499]=32'h10800040; 
ram[2500]=32'h00000000; 
ram[2501]=32'h27bdffc8; 
ram[2502]=32'hafbf0034; 
ram[2503]=32'hafb10030; 
ram[2504]=32'hafb0002c; 
ram[2505]=32'h04800036; 
ram[2506]=32'h00000000; 
ram[2507]=32'h00004821; 
ram[2508]=32'h3c056666; 
ram[2509]=32'h00003021; 
ram[2510]=32'h24a56667; 
ram[2511]=32'h0bc009d2; 
ram[2512]=32'h00000000; 
ram[2513]=32'h02003021; 
ram[2514]=32'h00850018; 
ram[2515]=32'h000417c3; 
ram[2516]=32'h00001810; 
ram[2517]=32'h00850018; 
ram[2518]=32'h00031883; 
ram[2519]=32'h00621823; 
ram[2520]=32'h00033840; 
ram[2521]=32'h00004010; 
ram[2522]=32'h000318c0; 
ram[2523]=32'h00e31821; 
ram[2524]=32'h00831823; 
ram[2525]=32'h24d00001; 
ram[2526]=32'h27a40018; 
ram[2527]=32'h00084083; 
ram[2528]=32'h00903821; 
ram[2529]=32'h24630030; 
ram[2530]=32'h01022023; 
ram[2531]=32'ha0e3ffff; 
ram[2532]=32'h1480ffec; 
ram[2533]=32'h00000000; 
ram[2534]=32'h15200012; 
ram[2535]=32'h00000000; 
ram[2536]=32'h2610ffff; 
ram[2537]=32'h2411ffff; 
ram[2538]=32'h27a40018; 
ram[2539]=32'h00901021; 
ram[2540]=32'h80440000; 
ram[2541]=32'h2610ffff; 
ram[2542]=32'h0fc00224; 
ram[2543]=32'h00000000; 
ram[2544]=32'h1611fff9; 
ram[2545]=32'h00000000; 
ram[2546]=32'h8fbf0034; 
ram[2547]=32'h8fb10030; 
ram[2548]=32'h8fb0002c; 
ram[2549]=32'h2404000a; 
ram[2550]=32'h27bd0038; 
ram[2551]=32'h0bc00224; 
ram[2552]=32'h00000000; 
ram[2553]=32'h27a30018; 
ram[2554]=32'h00701021; 
ram[2555]=32'h2403002d; 
ram[2556]=32'h24d00002; 
ram[2557]=32'ha0430000; 
ram[2558]=32'h0bc009e8; 
ram[2559]=32'h00000000; 
ram[2560]=32'h00042023; 
ram[2561]=32'h24090001; 
ram[2562]=32'h0bc009cc; 
ram[2563]=32'h00000000; 
ram[2564]=32'h24040030; 
ram[2565]=32'h0bc00224; 
ram[2566]=32'h00000000; 
ram[2567]=32'h27bdffd0; 
ram[2568]=32'h27a20018; 
ram[2569]=32'h3c059f00; 
ram[2570]=32'h27a60020; 
ram[2571]=32'hafb10028; 
ram[2572]=32'hafbf002c; 
ram[2573]=32'hafb00024; 
ram[2574]=32'h00408821; 
ram[2575]=32'h24a52920; 
ram[2576]=32'h3083000f; 
ram[2577]=32'h00a31821; 
ram[2578]=32'h90630000; 
ram[2579]=32'h24420001; 
ram[2580]=32'ha043ffff; 
ram[2581]=32'h00042102; 
ram[2582]=32'h1446fff9; 
ram[2583]=32'h00000000; 
ram[2584]=32'h27b0001f; 
ram[2585]=32'h2631ffff; 
ram[2586]=32'h82040000; 
ram[2587]=32'h2610ffff; 
ram[2588]=32'h0fc00224; 
ram[2589]=32'h00000000; 
ram[2590]=32'h1611fffb; 
ram[2591]=32'h00000000; 
ram[2592]=32'h8fbf002c; 
ram[2593]=32'h8fb10028; 
ram[2594]=32'h8fb00024; 
ram[2595]=32'h2404000a; 
ram[2596]=32'h27bd0030; 
ram[2597]=32'h0bc00224; 
ram[2598]=32'h00000000; 
ram[2599]=32'h00000000; 
ram[2600]=32'h72646461; 
ram[2601]=32'h25783020; 
ram[2602]=32'h78253d78; 
ram[2603]=32'h0000000a; 
ram[2604]=32'h65707974; 
ram[2605]=32'h6365723a; 
ram[2606]=32'h65766965; 
ram[2607]=32'h6e696220; 
ram[2608]=32'h6c696620; 
ram[2609]=32'h000a2e65; 
ram[2610]=32'h676e656c; 
ram[2611]=32'h3d206874; 
ram[2612]=32'h0a782520; 
ram[2613]=32'h00000000; 
ram[2614]=32'h72646461; 
ram[2615]=32'h25203d20; 
ram[2616]=32'h00000a78; 
ram[2617]=32'h65707974; 
ram[2618]=32'h6f6f623a; 
ram[2619]=32'h000a2074; 
ram[2620]=32'h6f746f67; 
ram[2621]=32'h64646120; 
ram[2622]=32'h203d2072; 
ram[2623]=32'h000a7825; 
ram[2624]=32'h200f3f3f; 
ram[2625]=32'h02040810; 
ram[2626]=32'he5e50001; 
ram[2627]=32'h0fffffff; 
ram[2628]=32'h0ffffff8; 
ram[2629]=32'h0fffffff; 
ram[2630]=32'hfffffff8; 
ram[2631]=32'h000055aa; 
ram[2632]=32'h33323130; 
ram[2633]=32'h37363534; 
ram[2634]=32'h62613938; 
ram[2635]=32'h66656463; 
ram[2636]=32'h33323130; 
ram[2637]=32'h37363534; 
ram[2638]=32'h42413938; 
ram[2639]=32'h46454443; 
ram[2640]=32'h00000000; 
ram[2641]=32'h00000000; 
ram[2642]=32'h00000000; 
ram[2643]=32'h00000000; 


	end
	
	reg[31:0] q;
	always_ff@(posedge clk_i)
	begin
	if(we_i) 
		begin
			if(be_i[0]) ram[adr_i][0] <= dat_i[7:0];
			if(be_i[1]) ram[adr_i][1] <= dat_i[15:8];
			if(be_i[2]) ram[adr_i][2] <= dat_i[23:16];
			if(be_i[3]) ram[adr_i][3] <= dat_i[31:24];
		end
		q <= ram[adr_i];
	end
	
	assign dat_o = q;
endmodule
