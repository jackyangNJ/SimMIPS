module const_base(
	output [31:0]base
);

	assign base = 32'd512;

endmodule