module SinglePortRam
(
	input clk_i,
	input we_i,
	input [11:0] adr_i, 
	input [3:0] be_i, 
	input [31:0] dat_i,
	output[31:0] dat_o
);
	
	// use a multi-dimensional packed array
	//to model individual bytes within the word
	// (* ram_init_file = "ram_init.mif" *) logic [3:0][7:0] ram[0:4095];
	logic [3:0][7:0] ram[0:4095];
	integer i;
	initial
	begin
		for(i=0;i<4096;i=i+1)
			ram[i] = 0;
ram[0]=32'h3c1d8000; 
ram[1]=32'h27bd13e0; 
ram[2]=32'h3c198000; 
ram[3]=32'h27390210; 
ram[4]=32'h0320f809; 
ram[5]=32'h1000ffff; 
ram[6]=32'h3c02b800; 
ram[7]=32'h2403ff80; 
ram[8]=32'ha04003f9; 
ram[9]=32'ha04303fb; 
ram[10]=32'h2403001b; 
ram[11]=32'ha04303f8; 
ram[12]=32'h24030003; 
ram[13]=32'ha04003f9; 
ram[14]=32'ha04303fb; 
ram[15]=32'h2403ffc7; 
ram[16]=32'ha04303fa; 
ram[17]=32'h2403000b; 
ram[18]=32'ha04303fc; 
ram[19]=32'h03e00008; 
ram[20]=32'h00000000; 
ram[21]=32'h308400ff; 
ram[22]=32'h3c02b800; 
ram[23]=32'h904303fd; 
ram[24]=32'h30630020; 
ram[25]=32'h1060fffc; 
ram[26]=32'h00000000; 
ram[27]=32'ha04403f8; 
ram[28]=32'h03e00008; 
ram[29]=32'h00000000; 
ram[30]=32'h90860000; 
ram[31]=32'h3c02b800; 
ram[32]=32'h10c0000a; 
ram[33]=32'h00000000; 
ram[34]=32'h904303fd; 
ram[35]=32'h30630020; 
ram[36]=32'h1060fffd; 
ram[37]=32'h00000000; 
ram[38]=32'ha04603f8; 
ram[39]=32'h24840001; 
ram[40]=32'h90860000; 
ram[41]=32'h14c0fff8; 
ram[42]=32'h00000000; 
ram[43]=32'h03e00008; 
ram[44]=32'h00000000; 
ram[45]=32'h3c02b800; 
ram[46]=32'h90420021; 
ram[47]=32'h304200ff; 
ram[48]=32'h03e00008; 
ram[49]=32'h00000000; 
ram[50]=32'h3c02b800; 
ram[51]=32'h2403000b; 
ram[52]=32'ha0430020; 
ram[53]=32'h90420020; 
ram[54]=32'h304200ff; 
ram[55]=32'h03e00008; 
ram[56]=32'h00000000; 
ram[57]=32'h3c02b800; 
ram[58]=32'h2403000a; 
ram[59]=32'ha0430020; 
ram[60]=32'h90420020; 
ram[61]=32'h304200ff; 
ram[62]=32'h03e00008; 
ram[63]=32'h00000000; 
ram[64]=32'h3c02b800; 
ram[65]=32'h2403000c; 
ram[66]=32'ha0430020; 
ram[67]=32'h90420020; 
ram[68]=32'h304200ff; 
ram[69]=32'h03e00008; 
ram[70]=32'h00000000; 
ram[71]=32'h3c02b800; 
ram[72]=32'h2403000c; 
ram[73]=32'ha04300a0; 
ram[74]=32'h904200a0; 
ram[75]=32'h304200ff; 
ram[76]=32'h03e00008; 
ram[77]=32'h00000000; 
ram[78]=32'h40026000; 
ram[79]=32'h3442ff00; 
ram[80]=32'h40826000; 
ram[81]=32'h3c02b800; 
ram[82]=32'h2408ffff; 
ram[83]=32'ha0480021; 
ram[84]=32'h2403000a; 
ram[85]=32'ha04800a1; 
ram[86]=32'h24070011; 
ram[87]=32'h24060002; 
ram[88]=32'h24050003; 
ram[89]=32'h24040068; 
ram[90]=32'h24080004; 
ram[91]=32'ha0470020; 
ram[92]=32'ha0460021; 
ram[93]=32'ha0480021; 
ram[94]=32'ha0450021; 
ram[95]=32'ha04700a0; 
ram[96]=32'ha04300a1; 
ram[97]=32'ha04600a1; 
ram[98]=32'ha04500a1; 
ram[99]=32'ha0440020; 
ram[100]=32'ha0430020; 
ram[101]=32'ha04400a0; 
ram[102]=32'ha04300a0; 
ram[103]=32'h03e00008; 
ram[104]=32'h00000000; 
ram[105]=32'h3c03b800; 
ram[106]=32'h2404000c; 
ram[107]=32'ha0640020; 
ram[108]=32'h90620020; 
ram[109]=32'h24050002; 
ram[110]=32'h30420007; 
ram[111]=32'h1045000e; 
ram[112]=32'h00000000; 
ram[113]=32'h24040007; 
ram[114]=32'h14440009; 
ram[115]=32'h00000000; 
ram[116]=32'h2404000b; 
ram[117]=32'ha0640020; 
ram[118]=32'h90640020; 
ram[119]=32'h2403ffff; 
ram[120]=32'h00042600; 
ram[121]=32'h00042603; 
ram[122]=32'h28840000; 
ram[123]=32'h0064100a; 
ram[124]=32'h03e00008; 
ram[125]=32'h00000000; 
ram[126]=32'ha06400a0; 
ram[127]=32'h906200a0; 
ram[128]=32'h30420007; 
ram[129]=32'h24420008; 
ram[130]=32'h03e00008; 
ram[131]=32'h00000000; 
ram[132]=32'h27bdffe0; 
ram[133]=32'hafbf001c; 
ram[134]=32'hafb20018; 
ram[135]=32'hafb10014; 
ram[136]=32'hafb00010; 
ram[137]=32'h0c000006; 
ram[138]=32'h00000000; 
ram[139]=32'h00001021; 
ram[140]=32'h40826000; 
ram[141]=32'h3c04ffff; 
ram[142]=32'h3c128000; 
ram[143]=32'h0c0000bc; 
ram[144]=32'h00000000; 
ram[145]=32'h00008021; 
ram[146]=32'h265203d8; 
ram[147]=32'h080000a0; 
ram[148]=32'h00000000; 
ram[149]=32'h0c000015; 
ram[150]=32'h00000000; 
ram[151]=32'h2404000a; 
ram[152]=32'h0c000015; 
ram[153]=32'h00000000; 
ram[154]=32'h26040010; 
ram[155]=32'h0c0000c2; 
ram[156]=32'h00000000; 
ram[157]=32'h26100001; 
ram[158]=32'h2a020010; 
ram[159]=32'h0002800a; 
ram[160]=32'h02002021; 
ram[161]=32'h0c0000d3; 
ram[162]=32'h00000000; 
ram[163]=32'h02402021; 
ram[164]=32'h00408821; 
ram[165]=32'h0c00001e; 
ram[166]=32'h00000000; 
ram[167]=32'h26040030; 
ram[168]=32'h308400ff; 
ram[169]=32'h0c000015; 
ram[170]=32'h00000000; 
ram[171]=32'h2404003d; 
ram[172]=32'h0c000015; 
ram[173]=32'h00000000; 
ram[174]=32'h24040031; 
ram[175]=32'h1620ffe5; 
ram[176]=32'h00000000; 
ram[177]=32'h24040030; 
ram[178]=32'h0c000015; 
ram[179]=32'h00000000; 
ram[180]=32'h2404000a; 
ram[181]=32'h0c000015; 
ram[182]=32'h00000000; 
ram[183]=32'h26040010; 
ram[184]=32'h0c0000ca; 
ram[185]=32'h00000000; 
ram[186]=32'h0800009d; 
ram[187]=32'h00000000; 
ram[188]=32'h3c02b800; 
ram[189]=32'h2403ffff; 
ram[190]=32'hac440404; 
ram[191]=32'hac430400; 
ram[192]=32'h03e00008; 
ram[193]=32'h00000000; 
ram[194]=32'h3c02b800; 
ram[195]=32'h8c430400; 
ram[196]=32'h24050001; 
ram[197]=32'h00852004; 
ram[198]=32'h00831825; 
ram[199]=32'hac430400; 
ram[200]=32'h03e00008; 
ram[201]=32'h00000000; 
ram[202]=32'h3c02b800; 
ram[203]=32'h24050001; 
ram[204]=32'h8c430400; 
ram[205]=32'h00852004; 
ram[206]=32'h00042827; 
ram[207]=32'h00a31824; 
ram[208]=32'hac430400; 
ram[209]=32'h03e00008; 
ram[210]=32'h00000000; 
ram[211]=32'h3c02b800; 
ram[212]=32'h8c430400; 
ram[213]=32'h24020001; 
ram[214]=32'h00821004; 
ram[215]=32'h00431024; 
ram[216]=32'h03e00008; 
ram[217]=32'h00000000; 
ram[218]=32'h27bdffe8; 
ram[219]=32'hafbf0014; 
ram[220]=32'h40046800; 
ram[221]=32'h0004202b; 
ram[222]=32'h0c000015; 
ram[223]=32'h00000000; 
ram[224]=32'h0c000040; 
ram[225]=32'h00000000; 
ram[226]=32'h00402021; 
ram[227]=32'h0c000015; 
ram[228]=32'h00000000; 
ram[229]=32'h3c02b800; 
ram[230]=32'h90440060; 
ram[231]=32'h8fbf0014; 
ram[232]=32'h308400ff; 
ram[233]=32'h27bd0018; 
ram[234]=32'h08000015; 
ram[235]=32'h00000000; 
ram[236]=32'h3c038000; 
ram[237]=32'h24630368; 
ram[238]=32'h00031900; 
ram[239]=32'h3c020800; 
ram[240]=32'h00031982; 
ram[241]=32'h00621825; 
ram[242]=32'h3c028000; 
ram[243]=32'hac430000; 
ram[244]=32'h03e00008; 
ram[245]=32'h00000000; 
ram[246]=32'h74726f70; 
ram[247]=32'h00000000; 

	end
	
	reg[31:0] q;
	always_ff@(posedge clk_i)
	begin
	if(we_i) 
		begin
			if(be_i[0]) ram[adr_i][0] <= dat_i[7:0];
			if(be_i[1]) ram[adr_i][1] <= dat_i[15:8];
			if(be_i[2]) ram[adr_i][2] <= dat_i[23:16];
			if(be_i[3]) ram[adr_i][3] <= dat_i[31:24];
		end
		q <= ram[adr_i];
	end
	
	assign dat_o = q;
endmodule
